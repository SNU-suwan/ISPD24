VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.69 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.127 0.078 0.525 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.114 0.334 0.64 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.114 0.162 0.27 0.19 ;
      RECT 0.242 0.162 0.27 0.428 ;
      RECT 0.114 0.162 0.142 0.544 ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X2 0 0 ;
  SIZE 0.448 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.262 0.083 0.506 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.512 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.078 0.338 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.082 0.166 0.27 0.194 ;
      RECT 0.242 0.166 0.27 0.602 ;
      RECT 0.054 0.574 0.27 0.602 ;
  END
END AND2_X2

MACRO AND3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X1 0 0 ;
  SIZE 0.512 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.173 0.192 0.211 0.568 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.192 0.08 0.576 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.576 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.114 0.462 0.654 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.274 0.105 0.398 0.137 ;
      RECT 0.37 0.105 0.398 0.664 ;
      RECT 0.054 0.636 0.398 0.664 ;
    LAYER M1 ;
      RECT 0.079 0.1 0.238 0.132 ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X2 0 0 ;
  SIZE 0.512 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.32 0.206 0.513 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.256 0.083 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.302 0.27 0.531 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.078 0.402 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.146 0.224 0.334 0.252 ;
      RECT 0.306 0.224 0.334 0.599 ;
      RECT 0.054 0.567 0.334 0.599 ;
    LAYER M1 ;
      RECT 0.048 0.078 0.08 0.188 ;
      RECT 0.048 0.156 0.298 0.188 ;
  END
END AND3_X2

MACRO AND4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_X1 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.576 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.114 0.526 0.654 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.192 0.272 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.142 0.512 ;
    END
  END A3
  OBS
    LAYER M1 ;
      RECT 0.141 0.104 0.298 0.152 ;
    LAYER M1 ;
      RECT 0.338 0.1 0.462 0.132 ;
      RECT 0.434 0.1 0.462 0.668 ;
      RECT 0.082 0.636 0.462 0.668 ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_X2 0 0 ;
  SIZE 0.64 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.577 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.241 0.398 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.192 0.27 0.577 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.142 0.577 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.096 0.526 0.64 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.142 0.104 0.298 0.136 ;
      RECT 0.342 0.165 0.462 0.197 ;
      RECT 0.434 0.165 0.462 0.664 ;
      RECT 0.082 0.632 0.462 0.664 ;
  END
END AND4_X2

MACRO ANTENNA
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ANTENNA 0 0 ;
  SIZE 0.192 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.078 0.08 0.256 ;
        RECT 0.048 0.512 0.08 0.69 ;
        RECT 0.048 0.228 0.142 0.256 ;
        RECT 0.114 0.228 0.142 0.54 ;
        RECT 0.048 0.512 0.142 0.54 ;
    END
  END I
END ANTENNA

MACRO AOI21_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X1 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.512 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.104 0.142 0.536 ;
        RECT 0.114 0.104 0.306 0.136 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.192 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.134 0.078 0.512 ;
    END
  END A2
  OBS
    LAYER M1 ;
      RECT 0.048 0.58 0.298 0.612 ;
      RECT 0.048 0.58 0.08 0.69 ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X2 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.302 0.398 0.448 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.166 0.206 0.599 ;
        RECT 0.077 0.166 0.43 0.194 ;
        RECT 0.434 0.507 0.462 0.599 ;
        RECT 0.178 0.571 0.462 0.599 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.23 0.27 0.512 ;
        RECT 0.242 0.23 0.531 0.258 ;
        RECT 0.493 0.23 0.531 0.448 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.142 0.448 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.048 0.55 0.08 0.677 ;
      RECT 0.498 0.516 0.526 0.677 ;
      RECT 0.048 0.643 0.526 0.677 ;
      RECT 0.146 0.102 0.535 0.13 ;
  END
END AOI21_X2

MACRO AOI22_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X1 0 0 ;
  SIZE 0.448 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.192 0.27 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.485 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.564 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.198 0.142 0.576 ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.141 0.102 0.334 0.13 ;
        RECT 0.306 0.102 0.334 0.58 ;
    END
  END ZN
  OBS
    LAYER M1 ;
      RECT 0.37 0.553 0.398 0.664 ;
      RECT 0.082 0.632 0.398 0.664 ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X2 0 0 ;
  SIZE 0.768 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.206 0.27 0.32 ;
        RECT 0.242 0.206 0.718 0.234 ;
        RECT 0.37 0.206 0.398 0.6 ;
        RECT 0.626 0.463 0.654 0.6 ;
        RECT 0.37 0.568 0.654 0.6 ;
        RECT 0.69 0.104 0.718 0.235 ;
        RECT 0.37 0.206 0.718 0.235 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.274 0.462 0.512 ;
        RECT 0.434 0.274 0.718 0.302 ;
        RECT 0.69 0.274 0.718 0.489 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.37 0.59 0.512 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.306 0.334 0.526 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.242 0.078 0.512 ;
    END
  END B2
  OBS
    LAYER M1 ;
      RECT 0.086 0.104 0.362 0.136 ;
    LAYER M1 ;
      RECT 0.626 0.078 0.654 0.17 ;
      RECT 0.406 0.138 0.654 0.17 ;
      RECT 0.69 0.557 0.718 0.672 ;
      RECT 0.077 0.644 0.718 0.672 ;
  END
END AOI22_X2

MACRO BUF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X1 0 0 ;
  SIZE 0.32 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.114 0.272 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.114 0.078 0.142 0.558 ;
  END
END BUF_X1

MACRO BUF_X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X12 0 0 ;
  SIZE 1.28 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.236 0.08 0.515 ;
        RECT 0.048 0.366 0.426 0.398 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.29 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.29 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.104 1.168 0.132 ;
        RECT 1.136 0.104 1.168 0.664 ;
        RECT 0.466 0.636 1.168 0.664 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.112 0.098 0.144 0.217 ;
      RECT 0.112 0.185 0.49 0.217 ;
      RECT 0.462 0.368 0.966 0.4 ;
      RECT 0.462 0.185 0.49 0.583 ;
      RECT 0.098 0.551 0.49 0.583 ;
      RECT 0.098 0.551 0.157 0.67 ;
  END
END BUF_X12

MACRO BUF_X16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X16 0 0 ;
  SIZE 1.664 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.232 0.078 0.512 ;
        RECT 0.05 0.368 0.554 0.4 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.102 1.552 0.13 ;
        RECT 1.52 0.102 1.552 0.66 ;
        RECT 0.594 0.632 1.552 0.66 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.114 0.141 0.142 0.235 ;
      RECT 0.114 0.203 0.618 0.235 ;
      RECT 0.59 0.366 1.454 0.398 ;
      RECT 0.59 0.203 0.618 0.488 ;
      RECT 0.114 0.456 0.618 0.488 ;
      RECT 0.114 0.456 0.142 0.643 ;
  END
END BUF_X16

MACRO BUF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X2 0 0 ;
  SIZE 0.32 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.267 0.078 0.512 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.078 0.206 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.048 0.129 0.08 0.22 ;
      RECT 0.048 0.192 0.142 0.22 ;
      RECT 0.114 0.192 0.142 0.584 ;
      RECT 0.048 0.556 0.142 0.584 ;
      RECT 0.048 0.556 0.08 0.664 ;
  END
END BUF_X2

MACRO BUF_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X4 0 0 ;
  SIZE 0.512 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.242 0.206 0.526 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.104 0.4 0.132 ;
        RECT 0.368 0.104 0.4 0.664 ;
        RECT 0.21 0.636 0.4 0.664 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.082 0.168 0.27 0.196 ;
      RECT 0.242 0.168 0.27 0.6 ;
      RECT 0.082 0.572 0.27 0.6 ;
  END
END BUF_X4

MACRO BUF_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X8 0 0 ;
  SIZE 0.896 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
        RECT 0.05 0.366 0.298 0.398 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.1 0.784 0.132 ;
        RECT 0.752 0.1 0.784 0.668 ;
        RECT 0.342 0.636 0.784 0.668 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.112 0.13 0.144 0.216 ;
      RECT 0.112 0.184 0.384 0.216 ;
      RECT 0.352 0.339 0.666 0.371 ;
      RECT 0.352 0.184 0.384 0.571 ;
      RECT 0.112 0.539 0.384 0.571 ;
      RECT 0.112 0.539 0.144 0.639 ;
  END
END BUF_X8

MACRO CLKBUF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X1 0 0 ;
  SIZE 0.32 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.114 0.272 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.114 0.078 0.142 0.523 ;
  END
END CLKBUF_X1

MACRO CLKBUF_X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X12 0 0 ;
  SIZE 1.28 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.238 0.08 0.53 ;
        RECT 0.048 0.336 0.426 0.368 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.29 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.29 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.104 1.168 0.132 ;
        RECT 1.136 0.104 1.168 0.664 ;
        RECT 0.466 0.636 1.168 0.664 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.043 0.168 0.494 0.196 ;
      RECT 0.462 0.168 0.494 0.346 ;
      RECT 0.462 0.314 0.998 0.346 ;
      RECT 0.462 0.168 0.49 0.578 ;
      RECT 0.114 0.55 0.49 0.578 ;
      RECT 0.114 0.55 0.142 0.67 ;
  END
END CLKBUF_X12

MACRO CLKBUF_X16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X16 0 0 ;
  SIZE 1.664 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.222 0.078 0.526 ;
        RECT 0.05 0.326 0.554 0.358 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.087 1.552 0.145 ;
        RECT 1.52 0.087 1.552 0.681 ;
        RECT 0.594 0.623 1.552 0.681 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.114 0.141 0.142 0.233 ;
      RECT 0.114 0.205 0.645 0.233 ;
      RECT 0.604 0.316 1.454 0.344 ;
      RECT 0.604 0.205 0.645 0.56 ;
      RECT 0.114 0.528 0.645 0.56 ;
      RECT 0.114 0.528 0.142 0.638 ;
  END
END CLKBUF_X16

MACRO CLKBUF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X2 0 0 ;
  SIZE 0.32 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.296 0.078 0.512 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.078 0.206 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.048 0.129 0.08 0.22 ;
      RECT 0.048 0.192 0.142 0.22 ;
      RECT 0.114 0.192 0.142 0.584 ;
      RECT 0.048 0.556 0.142 0.584 ;
      RECT 0.048 0.556 0.08 0.664 ;
  END
END CLKBUF_X2

MACRO CLKBUF_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X4 0 0 ;
  SIZE 0.512 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.142 0.526 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.104 0.4 0.132 ;
        RECT 0.368 0.104 0.4 0.664 ;
        RECT 0.205 0.636 0.4 0.664 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.041 0.168 0.206 0.196 ;
      RECT 0.178 0.168 0.206 0.6 ;
      RECT 0.082 0.572 0.206 0.6 ;
  END
END CLKBUF_X4

MACRO CLKBUF_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X8 0 0 ;
  SIZE 0.896 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
        RECT 0.05 0.256 0.079 0.356 ;
        RECT 0.05 0.328 0.318 0.356 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.104 0.782 0.136 ;
        RECT 0.754 0.104 0.782 0.664 ;
        RECT 0.338 0.632 0.782 0.664 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.05 0.172 0.434 0.2 ;
      RECT 0.406 0.37 0.718 0.402 ;
      RECT 0.406 0.172 0.434 0.482 ;
      RECT 0.114 0.45 0.434 0.482 ;
      RECT 0.114 0.45 0.142 0.542 ;
  END
END CLKBUF_X8

MACRO CLKGATETST_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATETST_X1 0 0 ;
  SIZE 1.088 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.69 0.238 0.718 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.01 0.104 1.038 0.654 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.32 0.078 0.664 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.098 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.098 0.028 ;
    END
  END VSS
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.142 0.672 ;
    END
  END E
  OBS
    LAYER V1 ;
      RECT 0.178 0.466 0.206 0.494 ;
      RECT 0.242 0.402 0.27 0.43 ;
      RECT 0.37 0.402 0.398 0.43 ;
      RECT 0.462 0.466 0.49 0.494 ;
      RECT 0.626 0.402 0.654 0.43 ;
      RECT 0.762 0.402 0.79 0.43 ;
      RECT 0.946 0.402 0.974 0.43 ;
    LAYER M1 ;
      RECT 0.178 0.166 0.302 0.194 ;
      RECT 0.178 0.166 0.206 0.662 ;
      RECT 0.178 0.63 0.366 0.662 ;
      RECT 0.306 0.307 0.334 0.574 ;
      RECT 0.558 0.184 0.59 0.574 ;
      RECT 0.306 0.546 0.59 0.574 ;
      RECT 0.434 0.104 0.91 0.132 ;
      RECT 0.434 0.104 0.462 0.334 ;
      RECT 0.882 0.104 0.91 0.662 ;
      RECT 0.466 0.63 0.91 0.662 ;
    LAYER M1 ;
      RECT 0.048 0.102 0.238 0.13 ;
      RECT 0.048 0.102 0.08 0.213 ;
      RECT 0.242 0.264 0.27 0.541 ;
      RECT 0.37 0.242 0.398 0.502 ;
      RECT 0.462 0.372 0.494 0.51 ;
      RECT 0.626 0.168 0.755 0.196 ;
      RECT 0.626 0.168 0.654 0.592 ;
      RECT 0.626 0.556 0.75 0.592 ;
      RECT 0.754 0.248 0.782 0.502 ;
      RECT 0.754 0.474 0.846 0.502 ;
      RECT 0.818 0.474 0.846 0.584 ;
      RECT 0.946 0.226 0.974 0.574 ;
    LAYER MINT1 ;
      RECT 0.146 0.466 0.522 0.494 ;
      RECT 0.73 0.402 1.006 0.43 ;
    LAYER MINT1 ;
      RECT 0.21 0.402 0.686 0.43 ;
  END
END CLKGATETST_X1

MACRO DFFRNQN_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRNQN_X1 0 0 ;
  SIZE 1.536 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.546 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.546 0.028 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.224 0.394 1.252 0.666 ;
        RECT 1.458 0.078 1.486 0.666 ;
        RECT 1.224 0.638 1.486 0.666 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.704 0.274 1.326 0.302 ;
    END
  END RN
  OBS
    LAYER V1 ;
      RECT 0.114 0.53 0.142 0.558 ;
      RECT 0.178 0.21 0.206 0.238 ;
      RECT 0.37 0.21 0.398 0.238 ;
      RECT 0.498 0.53 0.526 0.558 ;
      RECT 0.53 0.21 0.558 0.238 ;
      RECT 0.736 0.274 0.764 0.302 ;
      RECT 0.946 0.53 0.974 0.558 ;
      RECT 1.074 0.53 1.102 0.558 ;
      RECT 1.074 0.21 1.102 0.238 ;
      RECT 1.266 0.274 1.294 0.302 ;
    LAYER M1 ;
      RECT 0.048 0.104 0.08 0.188 ;
      RECT 0.048 0.16 0.142 0.188 ;
      RECT 0.114 0.16 0.142 0.606 ;
      RECT 0.048 0.567 0.142 0.606 ;
      RECT 0.048 0.567 0.08 0.664 ;
      RECT 0.37 0.194 0.398 0.494 ;
      RECT 0.498 0.402 0.526 0.574 ;
      RECT 0.526 0.194 0.558 0.294 ;
      RECT 0.736 0.258 0.764 0.438 ;
      RECT 0.946 0.274 0.974 0.578 ;
      RECT 1.074 0.446 1.102 0.622 ;
      RECT 1.074 0.174 1.102 0.317 ;
      RECT 1.156 0.166 1.188 0.664 ;
      RECT 1.266 0.174 1.294 0.318 ;
    LAYER M1 ;
      RECT 0.178 0.078 0.206 0.69 ;
      RECT 0.306 0.078 0.334 0.69 ;
      RECT 0.53 0.632 0.814 0.672 ;
      RECT 0.434 0.102 0.828 0.13 ;
      RECT 0.8 0.102 0.828 0.438 ;
      RECT 0.434 0.102 0.462 0.67 ;
      RECT 0.576 0.33 0.604 0.534 ;
      RECT 0.576 0.506 0.91 0.534 ;
      RECT 0.882 0.078 0.91 0.672 ;
      RECT 1.01 0.102 1.363 0.13 ;
      RECT 1.335 0.102 1.363 0.366 ;
      RECT 1.01 0.102 1.038 0.67 ;
    LAYER MINT1 ;
      RECT 0.082 0.53 1.134 0.558 ;
      RECT 0.146 0.21 1.134 0.238 ;
  END
END DFFRNQN_X1

MACRO DFFRNQQN_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRNQQN_X1 0 0 ;
  SIZE 1.664 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.078 1.616 0.689 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.224 0.394 1.252 0.666 ;
        RECT 1.458 0.078 1.486 0.666 ;
        RECT 1.224 0.638 1.486 0.666 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.704 0.274 1.326 0.302 ;
    END
  END RN
  OBS
    LAYER V1 ;
      RECT 0.114 0.53 0.142 0.558 ;
      RECT 0.178 0.21 0.206 0.238 ;
      RECT 0.37 0.21 0.398 0.238 ;
      RECT 0.498 0.53 0.526 0.558 ;
      RECT 0.53 0.21 0.558 0.238 ;
      RECT 0.736 0.274 0.764 0.302 ;
      RECT 0.946 0.53 0.974 0.558 ;
      RECT 1.074 0.53 1.102 0.558 ;
      RECT 1.074 0.21 1.102 0.238 ;
      RECT 1.266 0.274 1.294 0.302 ;
    LAYER M1 ;
      RECT 0.048 0.104 0.08 0.188 ;
      RECT 0.048 0.16 0.142 0.188 ;
      RECT 0.114 0.16 0.142 0.606 ;
      RECT 0.048 0.567 0.142 0.606 ;
      RECT 0.048 0.567 0.08 0.664 ;
      RECT 0.37 0.194 0.398 0.494 ;
      RECT 0.498 0.402 0.526 0.574 ;
      RECT 0.526 0.194 0.558 0.294 ;
      RECT 0.736 0.258 0.764 0.438 ;
      RECT 0.946 0.274 0.974 0.578 ;
      RECT 1.074 0.446 1.102 0.622 ;
      RECT 1.074 0.174 1.102 0.317 ;
      RECT 1.156 0.166 1.188 0.664 ;
      RECT 1.266 0.174 1.294 0.318 ;
    LAYER M1 ;
      RECT 0.178 0.078 0.206 0.69 ;
      RECT 0.306 0.078 0.334 0.69 ;
      RECT 0.53 0.632 0.814 0.672 ;
      RECT 0.434 0.102 0.828 0.13 ;
      RECT 0.8 0.102 0.828 0.438 ;
      RECT 0.434 0.102 0.462 0.67 ;
      RECT 0.576 0.33 0.604 0.534 ;
      RECT 0.576 0.506 0.91 0.534 ;
      RECT 0.882 0.078 0.91 0.672 ;
      RECT 1.01 0.102 1.363 0.13 ;
      RECT 1.335 0.102 1.363 0.366 ;
      RECT 1.01 0.102 1.038 0.67 ;
    LAYER MINT1 ;
      RECT 0.082 0.53 1.134 0.558 ;
      RECT 0.146 0.21 1.134 0.238 ;
  END
END DFFRNQQN_X1

MACRO DFFRNQ_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRNQ_X1 0 0 ;
  SIZE 1.664 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.078 1.616 0.689 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.704 0.274 1.326 0.302 ;
    END
  END RN
  OBS
    LAYER V1 ;
      RECT 0.114 0.53 0.142 0.558 ;
      RECT 0.178 0.21 0.206 0.238 ;
      RECT 0.37 0.21 0.398 0.238 ;
      RECT 0.498 0.53 0.526 0.558 ;
      RECT 0.53 0.21 0.558 0.238 ;
      RECT 0.736 0.274 0.764 0.302 ;
      RECT 0.946 0.53 0.974 0.558 ;
      RECT 1.074 0.53 1.102 0.558 ;
      RECT 1.074 0.21 1.102 0.238 ;
      RECT 1.266 0.274 1.294 0.302 ;
    LAYER M1 ;
      RECT 0.048 0.104 0.08 0.188 ;
      RECT 0.048 0.16 0.142 0.188 ;
      RECT 0.114 0.16 0.142 0.606 ;
      RECT 0.048 0.567 0.142 0.606 ;
      RECT 0.048 0.567 0.08 0.664 ;
      RECT 0.37 0.194 0.398 0.494 ;
      RECT 0.498 0.402 0.526 0.574 ;
      RECT 0.526 0.194 0.558 0.294 ;
      RECT 0.736 0.258 0.764 0.438 ;
      RECT 0.946 0.274 0.974 0.578 ;
      RECT 1.074 0.446 1.102 0.622 ;
      RECT 1.074 0.174 1.102 0.317 ;
      RECT 1.156 0.166 1.188 0.664 ;
      RECT 1.266 0.174 1.294 0.318 ;
    LAYER M1 ;
      RECT 0.178 0.078 0.206 0.69 ;
      RECT 0.306 0.078 0.334 0.69 ;
      RECT 0.53 0.632 0.814 0.672 ;
      RECT 0.434 0.102 0.828 0.13 ;
      RECT 0.8 0.102 0.828 0.438 ;
      RECT 0.434 0.102 0.462 0.67 ;
      RECT 0.576 0.33 0.604 0.534 ;
      RECT 0.576 0.506 0.91 0.534 ;
      RECT 0.882 0.078 0.91 0.672 ;
      RECT 1.01 0.102 1.363 0.13 ;
      RECT 1.335 0.102 1.363 0.366 ;
      RECT 1.01 0.102 1.038 0.67 ;
      RECT 1.224 0.394 1.252 0.666 ;
      RECT 1.458 0.078 1.486 0.666 ;
      RECT 1.224 0.638 1.486 0.666 ;
    LAYER MINT1 ;
      RECT 0.082 0.53 1.134 0.558 ;
      RECT 0.146 0.21 1.134 0.238 ;
  END
END DFFRNQ_X1

MACRO DFFSNQN_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSNQN_X1 0 0 ;
  SIZE 1.536 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.546 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.546 0.028 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.202 0.394 1.23 0.6 ;
        RECT 1.458 0.078 1.486 0.6 ;
        RECT 1.202 0.572 1.486 0.6 ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.722 0.274 1.326 0.302 ;
    END
  END SN
  OBS
    LAYER V1 ;
      RECT 0.114 0.53 0.142 0.558 ;
      RECT 0.178 0.21 0.206 0.238 ;
      RECT 0.37 0.21 0.398 0.238 ;
      RECT 0.498 0.53 0.526 0.558 ;
      RECT 0.526 0.21 0.554 0.238 ;
      RECT 0.754 0.274 0.782 0.302 ;
      RECT 0.946 0.53 0.974 0.558 ;
      RECT 1.074 0.53 1.102 0.558 ;
      RECT 1.074 0.21 1.102 0.238 ;
      RECT 1.266 0.274 1.294 0.302 ;
    LAYER M1 ;
      RECT 0.045 0.104 0.083 0.199 ;
      RECT 0.045 0.16 0.142 0.199 ;
      RECT 0.114 0.16 0.142 0.606 ;
      RECT 0.048 0.567 0.142 0.606 ;
      RECT 0.048 0.567 0.08 0.664 ;
      RECT 0.37 0.194 0.398 0.494 ;
      RECT 0.498 0.402 0.526 0.59 ;
      RECT 0.526 0.194 0.554 0.305 ;
      RECT 0.754 0.258 0.782 0.366 ;
      RECT 0.608 0.274 0.636 0.602 ;
      RECT 0.608 0.574 0.91 0.602 ;
      RECT 0.882 0.104 0.91 0.664 ;
      RECT 0.878 0.574 0.91 0.664 ;
      RECT 1.01 0.114 1.38 0.142 ;
      RECT 1.352 0.114 1.38 0.366 ;
      RECT 1.01 0.114 1.038 0.664 ;
      RECT 1.106 0.636 1.39 0.664 ;
    LAYER M1 ;
      RECT 0.178 0.078 0.206 0.69 ;
      RECT 0.306 0.078 0.334 0.69 ;
      RECT 0.434 0.122 0.846 0.15 ;
      RECT 0.818 0.122 0.846 0.366 ;
      RECT 0.434 0.122 0.462 0.67 ;
      RECT 0.946 0.274 0.974 0.574 ;
      RECT 1.074 0.393 1.106 0.594 ;
      RECT 1.074 0.194 1.106 0.325 ;
      RECT 1.266 0.186 1.294 0.318 ;
    LAYER MINT1 ;
      RECT 0.082 0.53 1.134 0.558 ;
      RECT 0.146 0.21 1.134 0.238 ;
  END
END DFFSNQN_X1

MACRO DFFSNQQN_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSNQQN_X1 0 0 ;
  SIZE 1.664 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.078 1.616 0.69 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.202 0.394 1.23 0.6 ;
        RECT 1.458 0.078 1.486 0.6 ;
        RECT 1.202 0.572 1.486 0.6 ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.722 0.274 1.326 0.302 ;
    END
  END SN
  OBS
    LAYER V1 ;
      RECT 0.114 0.53 0.142 0.558 ;
      RECT 0.178 0.21 0.206 0.238 ;
      RECT 0.37 0.21 0.398 0.238 ;
      RECT 0.498 0.53 0.526 0.558 ;
      RECT 0.526 0.21 0.554 0.238 ;
      RECT 0.754 0.274 0.782 0.302 ;
      RECT 0.946 0.53 0.974 0.558 ;
      RECT 1.074 0.53 1.102 0.558 ;
      RECT 1.074 0.21 1.102 0.238 ;
      RECT 1.266 0.274 1.294 0.302 ;
    LAYER M1 ;
      RECT 0.045 0.104 0.083 0.199 ;
      RECT 0.045 0.16 0.142 0.199 ;
      RECT 0.114 0.16 0.142 0.606 ;
      RECT 0.048 0.567 0.142 0.606 ;
      RECT 0.048 0.567 0.08 0.664 ;
      RECT 0.37 0.194 0.398 0.494 ;
      RECT 0.498 0.402 0.526 0.59 ;
      RECT 0.526 0.194 0.554 0.305 ;
      RECT 0.754 0.258 0.782 0.366 ;
      RECT 0.608 0.274 0.636 0.602 ;
      RECT 0.608 0.574 0.91 0.602 ;
      RECT 0.882 0.104 0.91 0.664 ;
      RECT 0.878 0.574 0.91 0.664 ;
      RECT 1.01 0.114 1.38 0.142 ;
      RECT 1.352 0.114 1.38 0.366 ;
      RECT 1.01 0.114 1.038 0.664 ;
      RECT 1.106 0.636 1.39 0.664 ;
    LAYER M1 ;
      RECT 0.178 0.078 0.206 0.69 ;
      RECT 0.306 0.078 0.334 0.69 ;
      RECT 0.434 0.122 0.846 0.15 ;
      RECT 0.818 0.122 0.846 0.366 ;
      RECT 0.434 0.122 0.462 0.67 ;
      RECT 0.946 0.274 0.974 0.574 ;
      RECT 1.074 0.393 1.106 0.594 ;
      RECT 1.074 0.194 1.106 0.325 ;
      RECT 1.266 0.186 1.294 0.318 ;
    LAYER MINT1 ;
      RECT 0.082 0.53 1.134 0.558 ;
      RECT 0.146 0.21 1.134 0.238 ;
  END
END DFFSNQQN_X1

MACRO DFFSNQ_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSNQ_X1 0 0 ;
  SIZE 1.664 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.078 1.616 0.69 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.722 0.274 1.326 0.302 ;
    END
  END SN
  OBS
    LAYER V1 ;
      RECT 0.114 0.53 0.142 0.558 ;
      RECT 0.178 0.21 0.206 0.238 ;
      RECT 0.37 0.21 0.398 0.238 ;
      RECT 0.498 0.53 0.526 0.558 ;
      RECT 0.526 0.21 0.554 0.238 ;
      RECT 0.754 0.274 0.782 0.302 ;
      RECT 0.946 0.53 0.974 0.558 ;
      RECT 1.074 0.53 1.102 0.558 ;
      RECT 1.074 0.21 1.102 0.238 ;
      RECT 1.266 0.274 1.294 0.302 ;
    LAYER M1 ;
      RECT 0.045 0.104 0.083 0.199 ;
      RECT 0.045 0.16 0.142 0.199 ;
      RECT 0.114 0.16 0.142 0.606 ;
      RECT 0.048 0.567 0.142 0.606 ;
      RECT 0.048 0.567 0.08 0.664 ;
      RECT 0.37 0.194 0.398 0.494 ;
      RECT 0.498 0.402 0.526 0.59 ;
      RECT 0.526 0.194 0.554 0.305 ;
      RECT 0.754 0.258 0.782 0.366 ;
      RECT 0.608 0.274 0.636 0.602 ;
      RECT 0.608 0.574 0.91 0.602 ;
      RECT 0.882 0.104 0.91 0.664 ;
      RECT 0.878 0.574 0.91 0.664 ;
      RECT 1.01 0.114 1.38 0.142 ;
      RECT 1.352 0.114 1.38 0.366 ;
      RECT 1.01 0.114 1.038 0.664 ;
      RECT 1.106 0.636 1.39 0.664 ;
    LAYER M1 ;
      RECT 0.178 0.078 0.206 0.69 ;
      RECT 0.306 0.078 0.334 0.69 ;
      RECT 0.434 0.122 0.846 0.15 ;
      RECT 0.818 0.122 0.846 0.366 ;
      RECT 0.434 0.122 0.462 0.67 ;
      RECT 0.946 0.274 0.974 0.574 ;
      RECT 1.074 0.393 1.106 0.594 ;
      RECT 1.074 0.194 1.106 0.325 ;
      RECT 1.266 0.186 1.294 0.318 ;
      RECT 1.202 0.394 1.23 0.6 ;
      RECT 1.458 0.078 1.486 0.6 ;
      RECT 1.202 0.572 1.486 0.6 ;
    LAYER MINT1 ;
      RECT 0.082 0.53 1.134 0.558 ;
      RECT 0.146 0.21 1.134 0.238 ;
  END
END DFFSNQ_X1

MACRO FA_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA_X1 0 0 ;
  SIZE 1.536 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.146 0.21 1.262 0.238 ;
      LAYER M1 ;
        RECT 1.202 0.178 1.23 0.366 ;
        RECT 0.578 0.194 0.61 0.362 ;
        RECT 0.178 0.194 0.206 0.59 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.21 0.466 1.102 0.494 ;
      LAYER M1 ;
        RECT 1.04 0.274 1.072 0.526 ;
        RECT 0.656 0.402 0.684 0.526 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.458 0.114 1.486 0.654 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.818 0.207 0.846 0.64 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.546 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.546 0.028 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.082 0.402 1.321 0.43 ;
      LAYER M1 ;
        RECT 1.261 0.402 1.289 0.59 ;
        RECT 0.103 0.338 0.142 0.462 ;
        RECT 0.027 0.338 0.142 0.366 ;
        RECT 0.027 0.178 0.065 0.366 ;
    END
  END A
  OBS
    LAYER V1 ;
      RECT 0.114 0.402 0.142 0.43 ;
      RECT 0.178 0.21 0.206 0.238 ;
      RECT 0.242 0.466 0.27 0.494 ;
      RECT 0.306 0.274 0.334 0.302 ;
      RECT 0.429 0.338 0.457 0.366 ;
      RECT 0.498 0.402 0.526 0.43 ;
      RECT 0.58 0.21 0.608 0.238 ;
      RECT 0.656 0.466 0.684 0.494 ;
      RECT 0.729 0.274 0.757 0.302 ;
      RECT 0.882 0.21 0.91 0.238 ;
      RECT 0.951 0.402 0.979 0.43 ;
      RECT 1.042 0.466 1.07 0.494 ;
      RECT 1.138 0.338 1.166 0.366 ;
      RECT 1.202 0.21 1.23 0.238 ;
      RECT 1.261 0.402 1.289 0.43 ;
      RECT 1.33 0.338 1.358 0.366 ;
    LAYER M1 ;
      RECT 0.306 0.104 0.334 0.664 ;
      RECT 0.498 0.274 0.526 0.507 ;
      RECT 0.949 0.274 0.981 0.494 ;
      RECT 0.846 0.104 1.084 0.136 ;
      RECT 1.33 0.274 1.358 0.526 ;
    LAYER M1 ;
      RECT 0.242 0.274 0.27 0.59 ;
      RECT 0.427 0.274 0.459 0.507 ;
      RECT 0.37 0.1 0.618 0.132 ;
      RECT 0.37 0.575 0.656 0.603 ;
      RECT 0.37 0.575 0.398 0.69 ;
      RECT 0.624 0.575 0.656 0.69 ;
      RECT 0.729 0.244 0.767 0.464 ;
      RECT 0.882 0.194 0.91 0.366 ;
      RECT 0.882 0.562 1.038 0.59 ;
      RECT 0.882 0.562 0.91 0.69 ;
      RECT 1.01 0.562 1.038 0.69 ;
      RECT 1.138 0.078 1.166 0.69 ;
    LAYER MINT1 ;
      RECT 0.397 0.338 1.39 0.366 ;
    LAYER MINT1 ;
      RECT 0.274 0.274 0.789 0.302 ;
  END
END FA_X1

MACRO FILLTIE
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLTIE 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
END FILLTIE

MACRO FILL_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL_X1 0 0 ;
  SIZE 0.128 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.138 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.138 0.028 ;
    END
  END VSS
END FILL_X1

MACRO FILL_X16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL_X16 0 0 ;
  SIZE 1.088 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.098 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.098 0.028 ;
    END
  END VSS
END FILL_X16

MACRO FILL_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL_X2 0 0 ;
  SIZE 0.192 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
END FILL_X2

MACRO FILL_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL_X4 0 0 ;
  SIZE 0.32 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
END FILL_X4

MACRO FILL_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL_X8 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
END FILL_X8

MACRO HA_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HA_X1 0 0 ;
  SIZE 0.832 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.274 0.27 0.584 ;
        RECT 0.434 0.274 0.462 0.584 ;
        RECT 0.242 0.556 0.462 0.584 ;
    END
  END A
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.754 0.18 0.782 0.638 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.842 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.842 0.028 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.512 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.082 0.078 0.638 ;
    END
  END CO
  OBS
    LAYER M1 ;
      RECT 0.114 0.166 0.37 0.198 ;
      RECT 0.114 0.166 0.142 0.664 ;
      RECT 0.566 0.274 0.596 0.664 ;
      RECT 0.114 0.636 0.596 0.664 ;
    LAYER M1 ;
      RECT 0.338 0.102 0.622 0.13 ;
      RECT 0.406 0.184 0.66 0.216 ;
      RECT 0.632 0.184 0.66 0.462 ;
      RECT 0.498 0.184 0.53 0.6 ;
  END
END HA_X1

MACRO INV_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X1 0 0 ;
  SIZE 0.192 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.114 0.142 0.64 ;
    END
  END ZN
END INV_X1

MACRO INV_X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X12 0 0 ;
  SIZE 0.896 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.142 0.576 ;
        RECT 0.114 0.368 0.686 0.396 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.102 0.851 0.13 ;
        RECT 0.813 0.102 0.851 0.668 ;
        RECT 0.054 0.636 0.851 0.668 ;
    END
  END ZN
END INV_X12

MACRO INV_X16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X16 0 0 ;
  SIZE 1.152 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.563 ;
        RECT 0.05 0.37 0.942 0.398 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.162 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.162 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.1 1.07 0.132 ;
        RECT 1.038 0.1 1.07 0.681 ;
        RECT 0.054 0.622 1.07 0.681 ;
    END
  END ZN
END INV_X16

MACRO INV_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X2 0 0 ;
  SIZE 0.256 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.13 0.142 0.576 ;
    END
  END ZN
END INV_X2

MACRO INV_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X4 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.256 0.08 0.512 ;
        RECT 0.048 0.368 0.238 0.396 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.142 0.334 0.2 ;
        RECT 0.306 0.142 0.334 0.626 ;
        RECT 0.059 0.568 0.334 0.626 ;
    END
  END ZN
END INV_X4

MACRO INV_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X8 0 0 ;
  SIZE 0.64 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.194 0.142 0.576 ;
        RECT 0.114 0.352 0.494 0.411 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.11 0.595 0.138 ;
        RECT 0.557 0.11 0.595 0.659 ;
        RECT 0.041 0.631 0.595 0.659 ;
    END
  END ZN
END INV_X8

MACRO LHQ_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LHQ_X1 0 0 ;
  SIZE 0.896 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.16 0.27 0.512 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.818 0.13 0.846 0.638 ;
    END
  END Q
  OBS
    LAYER M1 ;
      RECT 0.178 0.142 0.206 0.584 ;
      RECT 0.306 0.46 0.34 0.584 ;
      RECT 0.178 0.556 0.34 0.584 ;
      RECT 0.388 0.114 0.494 0.173 ;
      RECT 0.466 0.114 0.494 0.664 ;
      RECT 0.754 0.306 0.782 0.664 ;
      RECT 0.274 0.636 0.782 0.664 ;
    LAYER M1 ;
      RECT 0.05 0.078 0.352 0.106 ;
      RECT 0.05 0.078 0.078 0.212 ;
      RECT 0.05 0.184 0.142 0.212 ;
      RECT 0.324 0.078 0.352 0.35 ;
      RECT 0.324 0.322 0.398 0.35 ;
      RECT 0.37 0.322 0.398 0.414 ;
      RECT 0.114 0.184 0.142 0.584 ;
      RECT 0.048 0.556 0.142 0.584 ;
      RECT 0.048 0.556 0.08 0.69 ;
      RECT 0.53 0.114 0.718 0.142 ;
      RECT 0.53 0.114 0.558 0.494 ;
      RECT 0.69 0.114 0.718 0.593 ;
  END
END LHQ_X1

MACRO MUX2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2_X1 0 0 ;
  SIZE 0.832 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.142 0.448 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.027 0.242 0.055 0.664 ;
        RECT 0.027 0.636 0.222 0.664 ;
      LAYER MINT1 ;
        RECT 0.118 0.636 0.394 0.664 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.842 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.842 0.028 ;
    END
  END VSS
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.242 0.59 0.526 ;
    END
  END I0
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.69 0.192 0.718 0.638 ;
    END
  END Z
  OBS
    LAYER V1 ;
      RECT 0.15 0.636 0.206 0.664 ;
      RECT 0.306 0.338 0.334 0.366 ;
      RECT 0.306 0.636 0.362 0.664 ;
      RECT 0.498 0.338 0.526 0.366 ;
    LAYER M1 ;
      RECT 0.498 0.274 0.526 0.428 ;
      RECT 0.37 0.104 0.782 0.132 ;
      RECT 0.754 0.104 0.782 0.494 ;
      RECT 0.37 0.104 0.398 0.6 ;
    LAYER M1 ;
      RECT 0.08 0.162 0.334 0.19 ;
      RECT 0.306 0.162 0.334 0.52 ;
      RECT 0.099 0.492 0.334 0.52 ;
      RECT 0.099 0.492 0.157 0.576 ;
      RECT 0.434 0.306 0.462 0.681 ;
      RECT 0.29 0.636 0.462 0.681 ;
    LAYER MINT1 ;
      RECT 0.274 0.338 0.558 0.366 ;
  END
END MUX2_X1

MACRO NAND2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X1 0 0 ;
  SIZE 0.256 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.574 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.574 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.133 0.142 0.638 ;
        RECT 0.176 0.078 0.208 0.192 ;
        RECT 0.114 0.133 0.208 0.192 ;
    END
  END ZN
END NAND2_X1

MACRO NAND2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X2 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.123 0.142 0.626 ;
        RECT 0.114 0.123 0.27 0.181 ;
        RECT 0.242 0.424 0.27 0.626 ;
        RECT 0.114 0.589 0.27 0.626 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.225 0.206 0.553 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.274 0.078 0.69 ;
        RECT 0.306 0.274 0.334 0.69 ;
        RECT 0.05 0.662 0.334 0.69 ;
    END
  END A2
END NAND2_X2

MACRO NAND3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X1 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.255 0.206 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.215 0.078 0.574 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.32 0.27 0.448 ;
    END
  END A1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.082 0.142 0.69 ;
        RECT 0.114 0.082 0.336 0.11 ;
        RECT 0.306 0.512 0.334 0.69 ;
        RECT 0.114 0.662 0.334 0.69 ;
        RECT 0.304 0.082 0.336 0.256 ;
    END
  END ZN
END NAND3_X1

MACRO NAND3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X2 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.186 0.462 0.626 ;
        RECT 0.027 0.568 0.494 0.626 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.32 0.526 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.301 0.253 0.339 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.142 0.512 ;
    END
  END A3
  OBS
    LAYER M1 ;
      RECT 0.05 0.177 0.366 0.209 ;
    LAYER M1 ;
      RECT 0.21 0.111 0.526 0.141 ;
      RECT 0.498 0.111 0.526 0.225 ;
  END
END NAND3_X2

MACRO NAND4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X1 0 0 ;
  SIZE 0.448 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.256 0.398 0.574 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.512 ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.574 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.448 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.512 0.142 0.69 ;
        RECT 0.306 0.164 0.334 0.69 ;
        RECT 0.114 0.631 0.334 0.69 ;
        RECT 0.365 0.078 0.403 0.192 ;
        RECT 0.306 0.164 0.403 0.192 ;
    END
  END ZN
END NAND4_X1

MACRO NAND4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X2 0 0 ;
  SIZE 0.704 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.261 0.078 0.516 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.555 0.144 0.664 ;
        RECT 0.434 0.294 0.462 0.576 ;
        RECT 0.434 0.548 0.59 0.576 ;
        RECT 0.562 0.548 0.59 0.664 ;
        RECT 0.112 0.636 0.59 0.664 ;
        RECT 0.434 0.294 0.654 0.322 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.358 0.594 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.34 0.398 0.526 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.242 0.206 0.512 ;
    END
  END A3
  OBS
    LAYER M1 ;
      RECT 0.146 0.166 0.494 0.194 ;
    LAYER M1 ;
      RECT 0.048 0.102 0.43 0.13 ;
      RECT 0.048 0.102 0.08 0.213 ;
      RECT 0.624 0.078 0.656 0.258 ;
      RECT 0.274 0.23 0.656 0.258 ;
  END
END NAND4_X2

MACRO NOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X1 0 0 ;
  SIZE 0.256 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.512 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.13 0.142 0.635 ;
        RECT 0.114 0.576 0.208 0.635 ;
        RECT 0.176 0.576 0.208 0.69 ;
    END
  END ZN
END NOR2_X1

MACRO NOR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X2 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.142 0.142 0.584 ;
        RECT 0.114 0.556 0.208 0.584 ;
        RECT 0.176 0.556 0.208 0.64 ;
        RECT 0.114 0.142 0.27 0.17 ;
        RECT 0.242 0.142 0.27 0.344 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.215 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.078 0.078 0.494 ;
        RECT 0.05 0.078 0.334 0.106 ;
        RECT 0.306 0.078 0.334 0.494 ;
    END
  END A2
END NOR2_X2

MACRO NOR3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X1 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.553 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.553 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.32 0.27 0.448 ;
    END
  END A1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.078 0.142 0.642 ;
        RECT 0.114 0.078 0.337 0.106 ;
        RECT 0.114 0.614 0.336 0.642 ;
        RECT 0.304 0.512 0.336 0.69 ;
        RECT 0.303 0.078 0.337 0.256 ;
    END
  END ZN
END NOR3_X1

MACRO NOR3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X2 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.163 0.462 0.576 ;
        RECT 0.086 0.163 0.49 0.203 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.256 0.526 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.513 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.519 ;
    END
  END A3
  OBS
    LAYER M1 ;
      RECT 0.086 0.558 0.38 0.59 ;
    LAYER M1 ;
      RECT 0.498 0.516 0.526 0.655 ;
      RECT 0.21 0.627 0.526 0.655 ;
  END
END NOR3_X2

MACRO NOR4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X1 0 0 ;
  SIZE 0.448 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.194 0.398 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.194 0.27 0.512 ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.574 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.574 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.078 0.144 0.162 ;
        RECT 0.112 0.078 0.334 0.108 ;
        RECT 0.306 0.078 0.334 0.604 ;
        RECT 0.306 0.576 0.403 0.604 ;
        RECT 0.365 0.576 0.403 0.69 ;
    END
  END ZN
END NOR4_X1

MACRO NOR4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X2 0 0 ;
  SIZE 0.704 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.256 0.594 0.404 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.242 0.398 0.438 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.516 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.102 0.144 0.213 ;
        RECT 0.434 0.192 0.462 0.468 ;
        RECT 0.112 0.102 0.59 0.13 ;
        RECT 0.562 0.102 0.59 0.22 ;
        RECT 0.434 0.192 0.59 0.22 ;
        RECT 0.434 0.44 0.663 0.468 ;
    END
  END ZN
  OBS
    LAYER M1 ;
      RECT 0.048 0.555 0.08 0.664 ;
      RECT 0.048 0.636 0.43 0.664 ;
      RECT 0.338 0.504 0.656 0.532 ;
      RECT 0.624 0.504 0.656 0.664 ;
    LAYER M1 ;
      RECT 0.21 0.568 0.494 0.6 ;
  END
END NOR4_X2

MACRO OAI21_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X1 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.634 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.576 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.142 0.668 ;
        RECT 0.114 0.636 0.298 0.668 ;
    END
  END ZN
  OBS
    LAYER M1 ;
      RECT 0.05 0.078 0.078 0.187 ;
      RECT 0.05 0.155 0.298 0.187 ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X2 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.365 0.32 0.403 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.53 ;
        RECT 0.498 0.283 0.526 0.53 ;
        RECT 0.242 0.502 0.526 0.53 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.142 0.525 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.168 0.206 0.6 ;
        RECT 0.029 0.568 0.426 0.6 ;
        RECT 0.178 0.168 0.462 0.196 ;
        RECT 0.434 0.168 0.462 0.283 ;
    END
  END ZN
  OBS
    LAYER M1 ;
      RECT 0.048 0.104 0.526 0.132 ;
      RECT 0.048 0.104 0.08 0.213 ;
      RECT 0.498 0.104 0.526 0.215 ;
      RECT 0.146 0.636 0.535 0.664 ;
  END
END OAI21_X2

MACRO OAI22_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X1 0 0 ;
  SIZE 0.448 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.192 0.206 0.512 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.182 0.334 0.664 ;
        RECT 0.141 0.636 0.334 0.664 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.199 0.27 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.279 0.398 0.576 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.192 0.08 0.576 ;
    END
  END B2
  OBS
    LAYER M1 ;
      RECT 0.05 0.101 0.398 0.131 ;
      RECT 0.37 0.101 0.398 0.211 ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X2 0 0 ;
  SIZE 0.768 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.142 0.512 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.386 0.27 0.558 ;
        RECT 0.37 0.168 0.398 0.558 ;
        RECT 0.37 0.168 0.654 0.2 ;
        RECT 0.626 0.168 0.654 0.305 ;
        RECT 0.242 0.53 0.718 0.558 ;
        RECT 0.69 0.53 0.718 0.664 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.256 0.462 0.494 ;
        RECT 0.69 0.279 0.718 0.494 ;
        RECT 0.434 0.466 0.718 0.494 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.256 0.59 0.398 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.242 0.334 0.486 ;
    END
  END B1
  OBS
    LAYER M1 ;
      RECT 0.086 0.625 0.362 0.657 ;
    LAYER M1 ;
      RECT 0.406 0.598 0.654 0.63 ;
      RECT 0.626 0.598 0.654 0.69 ;
      RECT 0.041 0.1 0.718 0.132 ;
      RECT 0.69 0.1 0.718 0.211 ;
  END
END OAI22_X2

MACRO OR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X1 0 0 ;
  SIZE 0.384 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.104 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.243 0.078 0.641 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.114 0.334 0.64 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.114 0.13 0.142 0.584 ;
      RECT 0.242 0.336 0.27 0.584 ;
      RECT 0.114 0.556 0.27 0.584 ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X2 0 0 ;
  SIZE 0.448 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.142 0.512 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.078 0.338 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.077 0.154 0.27 0.188 ;
      RECT 0.242 0.154 0.27 0.608 ;
      RECT 0.146 0.58 0.27 0.608 ;
  END
END OR2_X2

MACRO OR3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X1 0 0 ;
  SIZE 0.512 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.576 ;
    END
  END A1
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.192 0.08 0.576 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.114 0.462 0.654 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.176 0.192 0.208 0.576 ;
    END
  END A2
  OBS
    LAYER M1 ;
      RECT 0.086 0.632 0.234 0.664 ;
    LAYER M1 ;
      RECT 0.054 0.109 0.398 0.137 ;
      RECT 0.37 0.109 0.398 0.673 ;
      RECT 0.278 0.631 0.398 0.673 ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X2 0 0 ;
  SIZE 0.512 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.526 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.255 0.142 0.448 ;
    END
  END A1
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.231 0.27 0.448 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.078 0.402 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.06 0.155 0.334 0.187 ;
      RECT 0.306 0.155 0.334 0.537 ;
      RECT 0.141 0.505 0.334 0.537 ;
    LAYER M1 ;
      RECT 0.05 0.573 0.302 0.603 ;
      RECT 0.05 0.573 0.078 0.686 ;
  END
END OR3_X2

MACRO OR4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4_X1 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.576 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.114 0.526 0.64 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.192 0.272 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.198 0.142 0.576 ;
    END
  END A3
  OBS
    LAYER M1 ;
      RECT 0.146 0.617 0.298 0.655 ;
    LAYER M1 ;
      RECT 0.054 0.102 0.462 0.13 ;
      RECT 0.434 0.102 0.462 0.662 ;
      RECT 0.338 0.63 0.462 0.662 ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4_X2 0 0 ;
  SIZE 0.64 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.213 0.27 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.213 0.142 0.576 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.53 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.191 0.078 0.576 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.496 0.128 0.528 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.054 0.104 0.46 0.136 ;
      RECT 0.432 0.104 0.46 0.624 ;
      RECT 0.342 0.568 0.46 0.624 ;
    LAYER M1 ;
      RECT 0.146 0.623 0.302 0.681 ;
  END
END OR4_X2

MACRO SDFFRNQ_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRNQ_X1 0 0 ;
  SIZE 1.92 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.276 0.078 0.534 ;
    END
  END CLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.372 0.334 0.6 ;
        RECT 0.562 0.314 0.59 0.6 ;
        RECT 0.306 0.572 0.59 0.6 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.93 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.93 0.028 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.363 0.526 0.528 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.078 1.872 0.69 ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.363 0.398 0.512 ;
    END
  END SI
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.965 0.338 1.598 0.366 ;
    END
  END RN
  OBS
    LAYER V1 ;
      RECT 0.114 0.274 0.142 0.302 ;
      RECT 0.178 0.53 0.206 0.558 ;
      RECT 0.69 0.53 0.718 0.558 ;
      RECT 0.754 0.402 0.782 0.43 ;
      RECT 0.818 0.274 0.846 0.302 ;
      RECT 0.997 0.338 1.025 0.366 ;
      RECT 1.065 0.402 1.093 0.43 ;
      RECT 1.202 0.274 1.23 0.302 ;
      RECT 1.266 0.53 1.294 0.558 ;
      RECT 1.394 0.274 1.422 0.302 ;
      RECT 1.538 0.338 1.566 0.366 ;
    LAYER M1 ;
      RECT 0.178 0.125 0.206 0.574 ;
      RECT 0.69 0.387 0.718 0.59 ;
      RECT 0.818 0.257 0.85 0.469 ;
      RECT 0.69 0.166 0.942 0.194 ;
      RECT 0.69 0.166 0.718 0.276 ;
      RECT 0.991 0.242 1.025 0.422 ;
      RECT 0.79 0.632 1.066 0.664 ;
      RECT 0.904 0.274 0.932 0.518 ;
      RECT 1.134 0.104 1.166 0.518 ;
      RECT 0.904 0.49 1.166 0.518 ;
      RECT 1.266 0.178 1.294 0.574 ;
      RECT 1.394 0.178 1.422 0.494 ;
      RECT 1.536 0.154 1.568 0.416 ;
    LAYER M1 ;
      RECT 0.045 0.096 0.083 0.232 ;
      RECT 0.045 0.204 0.142 0.232 ;
      RECT 0.114 0.204 0.142 0.632 ;
      RECT 0.045 0.604 0.142 0.632 ;
      RECT 0.045 0.604 0.083 0.688 ;
      RECT 0.242 0.267 0.515 0.295 ;
      RECT 0.242 0.096 0.27 0.672 ;
      RECT 0.338 0.184 0.654 0.212 ;
      RECT 0.626 0.184 0.654 0.276 ;
      RECT 0.392 0.636 0.754 0.668 ;
      RECT 0.754 0.247 0.782 0.546 ;
      RECT 0.466 0.102 0.878 0.13 ;
      RECT 1.063 0.24 1.095 0.446 ;
      RECT 1.202 0.171 1.23 0.511 ;
      RECT 1.458 0.146 1.49 0.69 ;
      RECT 1.33 0.078 1.635 0.106 ;
      RECT 1.607 0.078 1.635 0.366 ;
      RECT 1.33 0.078 1.358 0.646 ;
      RECT 1.165 0.618 1.358 0.646 ;
      RECT 1.554 0.46 1.582 0.672 ;
      RECT 1.714 0.078 1.742 0.672 ;
      RECT 1.554 0.632 1.742 0.672 ;
    LAYER MINT1 ;
      RECT 0.722 0.402 1.125 0.43 ;
      RECT 0.082 0.274 1.454 0.302 ;
    LAYER MINT1 ;
      RECT 0.146 0.53 1.326 0.558 ;
  END
END SDFFRNQ_X1

MACRO SDFFSNQ_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSNQ_X1 0 0 ;
  SIZE 1.92 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.272 0.078 0.512 ;
    END
  END CLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.372 0.334 0.6 ;
        RECT 0.562 0.314 0.59 0.6 ;
        RECT 0.306 0.572 0.59 0.6 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.93 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.93 0.028 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.384 0.526 0.528 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.078 1.872 0.69 ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.363 0.398 0.512 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MINT1 ;
        RECT 0.958 0.338 1.586 0.366 ;
    END
  END SN
  OBS
    LAYER V1 ;
      RECT 0.114 0.274 0.142 0.302 ;
      RECT 0.178 0.53 0.206 0.558 ;
      RECT 0.654 0.53 0.682 0.558 ;
      RECT 0.754 0.402 0.782 0.43 ;
      RECT 0.834 0.274 0.862 0.302 ;
      RECT 0.99 0.338 1.018 0.366 ;
      RECT 1.059 0.402 1.087 0.43 ;
      RECT 1.202 0.274 1.23 0.302 ;
      RECT 1.266 0.53 1.294 0.558 ;
      RECT 1.394 0.274 1.422 0.302 ;
      RECT 1.526 0.338 1.554 0.366 ;
    LAYER M1 ;
      RECT 0.178 0.104 0.206 0.619 ;
      RECT 0.654 0.387 0.682 0.574 ;
      RECT 0.83 0.257 0.862 0.469 ;
      RECT 0.69 0.166 0.942 0.194 ;
      RECT 0.69 0.166 0.718 0.276 ;
      RECT 1.057 0.24 1.089 0.446 ;
      RECT 1.202 0.171 1.23 0.383 ;
      RECT 1.33 0.104 1.645 0.132 ;
      RECT 1.607 0.104 1.645 0.366 ;
      RECT 1.33 0.104 1.358 0.646 ;
      RECT 1.165 0.618 1.358 0.646 ;
      RECT 1.462 0.402 1.49 0.602 ;
      RECT 1.714 0.104 1.742 0.602 ;
      RECT 1.462 0.574 1.742 0.602 ;
    LAYER M1 ;
      RECT 0.048 0.078 0.08 0.228 ;
      RECT 0.048 0.2 0.142 0.228 ;
      RECT 0.114 0.2 0.142 0.632 ;
      RECT 0.048 0.604 0.142 0.632 ;
      RECT 0.048 0.604 0.08 0.688 ;
      RECT 0.242 0.266 0.51 0.295 ;
      RECT 0.434 0.266 0.51 0.296 ;
      RECT 0.242 0.082 0.27 0.686 ;
      RECT 0.338 0.184 0.654 0.212 ;
      RECT 0.626 0.184 0.654 0.276 ;
      RECT 0.392 0.636 0.746 0.668 ;
      RECT 0.754 0.238 0.782 0.547 ;
      RECT 0.466 0.102 0.878 0.13 ;
      RECT 0.98 0.322 1.018 0.419 ;
      RECT 0.898 0.274 0.926 0.515 ;
      RECT 1.138 0.098 1.166 0.515 ;
      RECT 0.898 0.487 1.166 0.515 ;
      RECT 1.008 0.487 1.04 0.69 ;
      RECT 1.266 0.178 1.294 0.574 ;
      RECT 1.394 0.178 1.422 0.402 ;
      RECT 1.526 0.184 1.554 0.403 ;
      RECT 1.402 0.638 1.646 0.666 ;
    LAYER MINT1 ;
      RECT 0.722 0.402 1.119 0.43 ;
      RECT 0.082 0.274 1.454 0.302 ;
    LAYER MINT1 ;
      RECT 0.146 0.53 1.326 0.558 ;
  END
END SDFFSNQ_X1

MACRO TBUF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X1 0 0 ;
  SIZE 0.704 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.142 0.52 ;
        RECT 0.242 0.306 0.27 0.52 ;
        RECT 0.114 0.492 0.27 0.52 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.37 0.462 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.078 0.656 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.274 0.166 0.398 0.194 ;
      RECT 0.37 0.166 0.398 0.664 ;
      RECT 0.56 0.376 0.588 0.664 ;
      RECT 0.146 0.636 0.588 0.664 ;
    LAYER M1 ;
      RECT 0.05 0.312 0.206 0.34 ;
      RECT 0.178 0.312 0.206 0.418 ;
      RECT 0.05 0.078 0.078 0.686 ;
      RECT 0.202 0.102 0.542 0.13 ;
      RECT 0.202 0.102 0.23 0.258 ;
      RECT 0.202 0.23 0.334 0.258 ;
      RECT 0.51 0.102 0.542 0.314 ;
      RECT 0.306 0.23 0.334 0.6 ;
      RECT 0.146 0.572 0.334 0.6 ;
  END
END TBUF_X1

MACRO TBUF_X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X12 0 0 ;
  SIZE 1.728 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.346 0.526 0.441 ;
        RECT 0.626 0.409 0.654 0.576 ;
        RECT 0.434 0.409 0.71 0.441 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.738 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.738 0.028 ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.142 0.538 ;
        RECT 0.242 0.306 0.27 0.538 ;
        RECT 0.114 0.51 0.27 0.538 ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.931 0.532 0.989 0.62 ;
        RECT 1.586 0.532 1.614 0.624 ;
        RECT 0.882 0.102 1.688 0.13 ;
        RECT 1.633 0.102 1.688 0.564 ;
        RECT 0.931 0.532 1.688 0.564 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.05 0.312 0.206 0.34 ;
      RECT 0.178 0.312 0.206 0.404 ;
      RECT 0.05 0.174 0.078 0.664 ;
      RECT 0.142 0.104 0.814 0.132 ;
      RECT 0.142 0.104 0.174 0.26 ;
      RECT 0.782 0.104 0.814 0.294 ;
      RECT 0.142 0.232 0.334 0.26 ;
      RECT 0.782 0.25 1.579 0.294 ;
      RECT 0.306 0.232 0.334 0.602 ;
      RECT 0.146 0.574 0.334 0.602 ;
    LAYER M1 ;
      RECT 0.274 0.168 0.398 0.196 ;
      RECT 0.783 0.378 1.557 0.426 ;
      RECT 0.37 0.168 0.398 0.666 ;
      RECT 0.783 0.356 0.839 0.666 ;
      RECT 0.146 0.638 0.839 0.666 ;
  END
END TBUF_X12

MACRO TBUF_X16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X16 0 0 ;
  SIZE 2.112 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.39 0.142 0.514 ;
        RECT 0.24 0.32 0.272 0.514 ;
        RECT 0.114 0.486 0.272 0.514 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.346 0.59 0.445 ;
        RECT 0.69 0.405 0.718 0.576 ;
        RECT 0.47 0.405 0.902 0.445 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 2.122 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 2.122 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.072 0.078 1.104 0.2 ;
        RECT 1.072 0.528 1.104 0.69 ;
        RECT 1.072 0.528 2.062 0.568 ;
        RECT 1.968 0.078 2 0.2 ;
        RECT 1.968 0.528 2 0.69 ;
        RECT 1.072 0.142 2.062 0.2 ;
        RECT 2.034 0.142 2.062 0.576 ;
        RECT 1.968 0.528 2.062 0.576 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.21 0.104 0.974 0.132 ;
      RECT 0.21 0.104 0.238 0.264 ;
      RECT 0.21 0.236 0.36 0.264 ;
      RECT 0.946 0.104 0.974 0.331 ;
      RECT 0.946 0.273 1.984 0.331 ;
      RECT 0.328 0.236 0.36 0.601 ;
      RECT 0.146 0.569 0.36 0.601 ;
    LAYER M1 ;
      RECT 0.05 0.262 0.174 0.29 ;
      RECT 0.142 0.262 0.174 0.346 ;
      RECT 0.05 0.078 0.078 0.6 ;
      RECT 0.274 0.168 0.426 0.2 ;
      RECT 0.946 0.412 1.966 0.452 ;
      RECT 0.398 0.168 0.426 0.666 ;
      RECT 0.946 0.412 0.974 0.666 ;
      RECT 0.146 0.638 0.974 0.666 ;
  END
END TBUF_X16

MACRO TBUF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X2 0 0 ;
  SIZE 0.768 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.142 0.532 ;
        RECT 0.242 0.306 0.27 0.532 ;
        RECT 0.114 0.504 0.27 0.532 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.382 0.462 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.078 0.656 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.274 0.166 0.398 0.194 ;
      RECT 0.37 0.166 0.398 0.664 ;
      RECT 0.498 0.443 0.53 0.664 ;
      RECT 0.146 0.636 0.53 0.664 ;
    LAYER M1 ;
      RECT 0.05 0.312 0.206 0.34 ;
      RECT 0.178 0.312 0.206 0.404 ;
      RECT 0.05 0.078 0.078 0.612 ;
      RECT 0.202 0.102 0.514 0.13 ;
      RECT 0.202 0.102 0.23 0.258 ;
      RECT 0.202 0.23 0.334 0.258 ;
      RECT 0.482 0.102 0.514 0.314 ;
      RECT 0.306 0.23 0.334 0.6 ;
      RECT 0.146 0.568 0.334 0.6 ;
  END
END TBUF_X2

MACRO TBUF_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X4 0 0 ;
  SIZE 0.96 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.346 0.462 0.594 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.97 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.97 0.028 ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.142 0.512 ;
        RECT 0.242 0.306 0.27 0.512 ;
        RECT 0.114 0.484 0.27 0.512 ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.688 0.078 0.72 0.256 ;
        RECT 0.688 0.524 0.72 0.69 ;
        RECT 0.688 0.524 0.91 0.552 ;
        RECT 0.816 0.524 0.848 0.69 ;
        RECT 0.813 0.078 0.851 0.256 ;
        RECT 0.688 0.224 0.91 0.256 ;
        RECT 0.882 0.224 0.91 0.583 ;
        RECT 0.816 0.524 0.91 0.583 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.05 0.312 0.206 0.34 ;
      RECT 0.178 0.312 0.206 0.404 ;
      RECT 0.05 0.104 0.078 0.594 ;
      RECT 0.202 0.104 0.574 0.132 ;
      RECT 0.202 0.104 0.23 0.26 ;
      RECT 0.202 0.232 0.334 0.26 ;
      RECT 0.534 0.292 0.838 0.32 ;
      RECT 0.534 0.104 0.574 0.348 ;
      RECT 0.306 0.232 0.334 0.602 ;
      RECT 0.146 0.568 0.334 0.602 ;
    LAYER M1 ;
      RECT 0.274 0.168 0.398 0.196 ;
      RECT 0.534 0.416 0.814 0.456 ;
      RECT 0.37 0.168 0.398 0.666 ;
      RECT 0.534 0.392 0.574 0.666 ;
      RECT 0.082 0.638 0.574 0.666 ;
  END
END TBUF_X4

MACRO TBUF_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X8 0 0 ;
  SIZE 1.344 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.142 0.512 ;
        RECT 0.306 0.32 0.334 0.512 ;
        RECT 0.114 0.484 0.334 0.512 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.354 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.354 0.028 ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.346 0.526 0.576 ;
        RECT 0.498 0.402 0.618 0.434 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.816 0.078 0.848 0.192 ;
        RECT 0.816 0.519 0.848 0.69 ;
        RECT 0.816 0.519 1.294 0.577 ;
        RECT 1.2 0.078 1.232 0.192 ;
        RECT 1.2 0.519 1.232 0.69 ;
        RECT 1.2 0.133 1.294 0.192 ;
        RECT 0.816 0.16 1.294 0.192 ;
        RECT 1.266 0.133 1.294 0.578 ;
        RECT 1.2 0.519 1.294 0.578 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.274 0.166 0.462 0.194 ;
      RECT 0.669 0.403 1.183 0.461 ;
      RECT 0.434 0.166 0.462 0.664 ;
      RECT 0.669 0.386 0.709 0.664 ;
      RECT 0.122 0.636 0.709 0.664 ;
    LAYER M1 ;
      RECT 0.05 0.312 0.23 0.34 ;
      RECT 0.186 0.312 0.23 0.43 ;
      RECT 0.05 0.078 0.078 0.638 ;
      RECT 0.2 0.102 0.718 0.13 ;
      RECT 0.2 0.102 0.232 0.258 ;
      RECT 0.2 0.23 0.398 0.258 ;
      RECT 0.69 0.258 1.198 0.286 ;
      RECT 0.69 0.102 0.718 0.342 ;
      RECT 0.37 0.23 0.398 0.6 ;
      RECT 0.146 0.572 0.398 0.6 ;
  END
END TBUF_X8

MACRO TIEH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEH 0 0 ;
  SIZE 0.192 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.473 0.147 0.69 ;
    END
  END Z
  OBS
    LAYER M1 ;
      RECT 0.114 0.104 0.142 0.429 ;
  END
END TIEH

MACRO TIEL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEL 0 0 ;
  SIZE 0.192 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.078 0.147 0.266 ;
    END
  END ZN
  OBS
    LAYER M1 ;
      RECT 0.114 0.336 0.142 0.664 ;
  END
END TIEL

MACRO XNOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_X1 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.248 0.462 0.59 ;
        RECT 0.274 0.558 0.462 0.59 ;
        RECT 0.302 0.166 0.531 0.194 ;
        RECT 0.493 0.166 0.531 0.276 ;
        RECT 0.434 0.248 0.531 0.276 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.252 0.206 0.432 ;
        RECT 0.178 0.252 0.398 0.28 ;
        RECT 0.37 0.252 0.398 0.432 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.242 0.078 0.69 ;
        RECT 0.498 0.32 0.526 0.69 ;
        RECT 0.05 0.662 0.526 0.69 ;
    END
  END A2
  OBS
    LAYER M1 ;
      RECT 0.114 0.184 0.234 0.216 ;
      RECT 0.246 0.34 0.274 0.496 ;
      RECT 0.114 0.468 0.274 0.496 ;
      RECT 0.114 0.184 0.142 0.556 ;
    LAYER M1 ;
      RECT 0.21 0.102 0.535 0.13 ;
  END
END XNOR2_X1

MACRO XOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_X1 0 0 ;
  SIZE 0.576 BY 0.768 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.274 0.177 0.462 0.209 ;
        RECT 0.434 0.177 0.462 0.52 ;
        RECT 0.434 0.492 0.528 0.52 ;
        RECT 0.496 0.492 0.528 0.602 ;
        RECT 0.315 0.574 0.528 0.602 ;
    END
  END Z
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.344 0.21 0.514 ;
        RECT 0.37 0.32 0.398 0.514 ;
        RECT 0.178 0.486 0.398 0.514 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.078 0.078 0.526 ;
        RECT 0.05 0.078 0.526 0.106 ;
        RECT 0.498 0.078 0.526 0.448 ;
    END
  END A2
  OBS
    LAYER M1 ;
      RECT 0.114 0.28 0.274 0.308 ;
      RECT 0.246 0.28 0.274 0.432 ;
      RECT 0.114 0.142 0.142 0.584 ;
      RECT 0.114 0.552 0.247 0.584 ;
    LAYER M1 ;
      RECT 0.246 0.638 0.535 0.666 ;
  END
END XOR2_X1

MACRO h3_mgc_des_perf_a
   CLASS BLOCK ;
   FOREIGN h3 ;
   ORIGIN 0 0 ;
   SIZE 175.744 BY 94.72 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1005_n_65753
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.434 0.163 24.462 ;
      END
   END FE_OFN1005_n_65753

   PIN FE_OFN1022_n_3701
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.33 0.163 9.358 ;
      END
   END FE_OFN1022_n_3701

   PIN FE_OFN1051_n_5643
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.938 0.163 77.966 ;
      END
   END FE_OFN1051_n_5643

   PIN FE_OFN106_n_95123
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.762 0.163 35.79 ;
      END
   END FE_OFN106_n_95123

   PIN FE_OFN1075_n_116
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.474 0.0 7.502 0.082 ;
      END
   END FE_OFN1075_n_116

   PIN FE_OFN1095_g303299_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.234 0.163 5.262 ;
      END
   END FE_OFN1095_g303299_p

   PIN FE_OFN1121_n_4882
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.002 0.163 78.03 ;
      END
   END FE_OFN1121_n_4882

   PIN FE_OFN1203_n_118585
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 57.01 0.0 57.038 0.082 ;
      END
   END FE_OFN1203_n_118585

   PIN FE_OFN1215_n_3935
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.298 0.163 5.326 ;
      END
   END FE_OFN1215_n_3935

   PIN FE_OFN1225_n_6583
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.738 0.0 26.766 0.163 ;
      END
   END FE_OFN1225_n_6583

   PIN FE_OFN1228_n_3045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.53 0.0 4.558 0.163 ;
      END
   END FE_OFN1228_n_3045

   PIN FE_OFN1431_n_22026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.914 0.0 12.942 0.163 ;
      END
   END FE_OFN1431_n_22026

   PIN FE_OFN1534_n_4068
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.362 0.163 5.39 ;
      END
   END FE_OFN1534_n_4068

   PIN FE_OFN1551_n_13938
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.482 0.163 10.51 ;
      END
   END FE_OFN1551_n_13938

   PIN FE_OFN1579_n_3047
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.426 0.163 5.454 ;
      END
   END FE_OFN1579_n_3047

   PIN FE_OFN1625_n_3863
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.49 0.163 5.518 ;
      END
   END FE_OFN1625_n_3863

   PIN FE_OFN1667_n_66371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.762 0.0 27.79 0.163 ;
      END
   END FE_OFN1667_n_66371

   PIN FE_OFN1863_n_4923
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.554 0.163 5.582 ;
      END
   END FE_OFN1863_n_4923

   PIN FE_OFN1930_n_18862
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.618 0.163 5.646 ;
      END
   END FE_OFN1930_n_18862

   PIN FE_OFN1959_n_6873
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.194 0.0 30.222 0.163 ;
      END
   END FE_OFN1959_n_6873

   PIN FE_OFN2010_n_27918
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.482 0.0 18.51 0.163 ;
      END
   END FE_OFN2010_n_27918

   PIN FE_OFN2014_n_23906
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.578 0.163 62.606 ;
      END
   END FE_OFN2014_n_23906

   PIN FE_OFN2148_n_118596
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.082 0.163 4.11 ;
      END
   END FE_OFN2148_n_118596

   PIN FE_OFN2171_n_117298
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.042 0.0 53.07 0.163 ;
      END
   END FE_OFN2171_n_117298

   PIN FE_OFN2175_n_21905
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.082 0.163 4.11 ;
      END
   END FE_OFN2175_n_21905

   PIN FE_OFN2254_n_23876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.146 0.163 4.174 ;
      END
   END FE_OFN2254_n_23876

   PIN FE_OFN2334_n_23919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.57 0.163 3.598 ;
      END
   END FE_OFN2334_n_23919

   PIN FE_OFN2352_n_27890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.138 0.0 33.166 0.163 ;
      END
   END FE_OFN2352_n_27890

   PIN FE_OFN2353_n_19056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.682 0.163 5.71 ;
      END
   END FE_OFN2353_n_19056

   PIN FE_OFN2395_n_61534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.746 0.163 5.774 ;
      END
   END FE_OFN2395_n_61534

   PIN FE_OFN2397_n_4104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.538 0.163 7.566 ;
      END
   END FE_OFN2397_n_4104

   PIN FE_OFN2400_n_18228
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.282 0.163 7.31 ;
      END
   END FE_OFN2400_n_18228

   PIN FE_OFN2418_n_26365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.882 0.0 16.91 0.163 ;
      END
   END FE_OFN2418_n_26365

   PIN FE_OFN2419_n_25888
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.09 0.163 55.118 ;
      END
   END FE_OFN2419_n_25888

   PIN FE_OFN2473_n_117820
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.714 0.0 105.742 0.163 ;
      END
   END FE_OFN2473_n_117820

   PIN FE_OFN2484_n_25794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.21 0.163 4.238 ;
      END
   END FE_OFN2484_n_25794

   PIN FE_OFN2502_n_5437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.266 0.0 25.294 0.163 ;
      END
   END FE_OFN2502_n_5437

   PIN FE_OFN2505_n_4918
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.642 0.163 62.67 ;
      END
   END FE_OFN2505_n_4918

   PIN FE_OFN2678_n_23958
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 81.778 0.163 81.806 ;
      END
   END FE_OFN2678_n_23958

   PIN FE_OFN2701_n_2549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.306 0.163 16.334 ;
      END
   END FE_OFN2701_n_2549

   PIN FE_OFN2720_n_25980
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.826 0.163 35.854 ;
      END
   END FE_OFN2720_n_25980

   PIN FE_OFN2787_n_5684
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.89 0.163 35.918 ;
      END
   END FE_OFN2787_n_5684

   PIN FE_OFN2790_n_4079
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.65 0.0 1.678 0.163 ;
      END
   END FE_OFN2790_n_4079

   PIN FE_OFN287_n_76853
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.858 0.0 7.886 0.163 ;
      END
   END FE_OFN287_n_76853

   PIN FE_OFN2929_n_4064
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.306 0.0 8.334 0.163 ;
      END
   END FE_OFN2929_n_4064

   PIN FE_OFN2976_n_65768
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.506 0.163 35.534 ;
      END
   END FE_OFN2976_n_65768

   PIN FE_OFN3004_n_4088
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.018 0.0 4.046 0.163 ;
      END
   END FE_OFN3004_n_4088

   PIN FE_OFN3018_n_69766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.97 0.0 97.998 0.163 ;
      END
   END FE_OFN3018_n_69766

   PIN FE_OFN3050_n_3016
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.146 0.163 20.174 ;
      END
   END FE_OFN3050_n_3016

   PIN FE_OFN3096_n_4811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.114 0.163 8.142 ;
      END
   END FE_OFN3096_n_4811

   PIN FE_OFN3163_n_2780
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.69 0.0 0.718 0.163 ;
      END
   END FE_OFN3163_n_2780

   PIN FE_OFN3206_n_32181
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.09 0.0 55.118 0.163 ;
      END
   END FE_OFN3206_n_32181

   PIN FE_OFN3230_n_3189
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.714 0.0 1.742 0.163 ;
      END
   END FE_OFN3230_n_3189

   PIN FE_OFN3235_n_2155
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.314 0.0 3.342 0.163 ;
      END
   END FE_OFN3235_n_2155

   PIN FE_OFN3241_n_4790
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.178 0.163 8.206 ;
      END
   END FE_OFN3241_n_4790

   PIN FE_OFN325_n_70684
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.322 0.0 94.35 0.163 ;
      END
   END FE_OFN325_n_70684

   PIN FE_OFN327_n_70685
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.938 0.0 101.966 0.163 ;
      END
   END FE_OFN327_n_70685

   PIN FE_OFN3364_n_25895
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.61 0.163 66.638 ;
      END
   END FE_OFN3364_n_25895

   PIN FE_OFN3366_n_5443
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 81.842 0.163 81.87 ;
      END
   END FE_OFN3366_n_5443

   PIN FE_OFN3464_n_67106
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.818 94.557 40.846 94.72 ;
      END
   END FE_OFN3464_n_67106

   PIN FE_OFN3486_n_1596
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.274 0.163 4.302 ;
      END
   END FE_OFN3486_n_1596

   PIN FE_OFN3517_n_23820
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.546 0.163 10.574 ;
      END
   END FE_OFN3517_n_23820

   PIN FE_OFN3531_n_19107
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.858 0.082 7.886 ;
      END
   END FE_OFN3531_n_19107

   PIN FE_OFN3549_n_7898
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.61 0.163 10.638 ;
      END
   END FE_OFN3549_n_7898

   PIN FE_OFN3617_n_18380
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.338 0.163 4.366 ;
      END
   END FE_OFN3617_n_18380

   PIN FE_OFN3628_n_4557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.274 0.163 28.302 ;
      END
   END FE_OFN3628_n_4557

   PIN FE_OFN3720_n_4799
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.634 0.163 3.662 ;
      END
   END FE_OFN3720_n_4799

   PIN FE_OFN3800_n_23840
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.81 0.163 5.838 ;
      END
   END FE_OFN3800_n_23840

   PIN FE_OFN3910_n_5532
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.066 0.163 78.094 ;
      END
   END FE_OFN3910_n_5532

   PIN FE_OFN4090_n_2663
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 5.746 0.163 5.774 ;
      END
   END FE_OFN4090_n_2663

   PIN FE_OFN4798_n_21953
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.874 0.163 5.902 ;
      END
   END FE_OFN4798_n_21953

   PIN FE_OFN666_n_31829
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.378 0.0 51.406 0.163 ;
      END
   END FE_OFN666_n_31829

   PIN FE_OFN693_n_27625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.058 0.0 11.086 0.163 ;
      END
   END FE_OFN693_n_27625

   PIN FE_OFN715_n_24030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.274 0.0 4.302 0.163 ;
      END
   END FE_OFN715_n_24030

   PIN FE_OFN737_n_4131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.938 0.163 5.966 ;
      END
   END FE_OFN737_n_4131

   PIN FE_OFN847_n_4294
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.002 0.163 6.03 ;
      END
   END FE_OFN847_n_4294

   PIN FE_OFN848_n_4958
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.37 0.163 16.398 ;
      END
   END FE_OFN848_n_4958

   PIN FE_OFN853_n_3353
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.066 0.163 6.094 ;
      END
   END FE_OFN853_n_3353

   PIN FE_OFN911_n_21872
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 5.81 0.163 5.838 ;
      END
   END FE_OFN911_n_21872

   PIN FE_OFN948_n_3795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.242 0.163 8.27 ;
      END
   END FE_OFN948_n_3795

   PIN FE_OFN965_n_25771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.13 0.163 6.158 ;
      END
   END FE_OFN965_n_25771

   PIN FE_OFN973_n_63299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.194 0.163 6.222 ;
      END
   END FE_OFN973_n_63299

   PIN FE_OFN975_n_2435
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.602 0.163 7.63 ;
      END
   END FE_OFN975_n_2435

   PIN g205805_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.226 0.0 74.254 0.163 ;
      END
   END g205805_da

   PIN g221053_u1_o
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.906 94.557 17.934 94.72 ;
      END
   END g221053_u1_o

   PIN g222840_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.674 0.163 10.702 ;
      END
   END g222840_p

   PIN g229165_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.45 0.0 102.478 0.163 ;
      END
   END g229165_p

   PIN g229250_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.514 0.0 102.542 0.163 ;
      END
   END g229250_p

   PIN g229781_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.41 0.0 23.438 0.163 ;
      END
   END g229781_p

   PIN g231281_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.21 0.163 20.238 ;
      END
   END g231281_p

   PIN g233246_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.506 0.0 11.534 0.163 ;
      END
   END g233246_p

   PIN g233290_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.498 0.163 16.526 ;
      END
   END g233290_p

   PIN g233318_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.202 0.0 25.23 0.163 ;
      END
   END g233318_p

   PIN g233379_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.986 0.0 24.014 0.163 ;
      END
   END g233379_p

   PIN g233525_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.794 0.163 39.822 ;
      END
   END g233525_p

   PIN g233666_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.53 0.163 12.558 ;
      END
   END g233666_p

   PIN g233787_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.074 0.163 9.102 ;
      END
   END g233787_p

   PIN g235027_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.698 0.0 19.726 0.163 ;
      END
   END g235027_p

   PIN g235236_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.234 0.0 21.262 0.163 ;
      END
   END g235236_p

   PIN g235278_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.89 0.0 19.918 0.163 ;
      END
   END g235278_p

   PIN g235292_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.01 0.0 25.038 0.163 ;
      END
   END g235292_p

   PIN g235499_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.154 0.163 55.182 ;
      END
   END g235499_p

   PIN g235503_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.506 0.0 19.534 0.163 ;
      END
   END g235503_p

   PIN g236596_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.186 0.0 11.214 0.163 ;
      END
   END g236596_da

   PIN g236596_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.33 0.0 9.358 0.163 ;
      END
   END g236596_db

   PIN g264946_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.706 0.0 86.734 0.163 ;
      END
   END g264946_da

   PIN g264946_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.962 0.0 86.99 0.163 ;
      END
   END g264946_db

   PIN g265666_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.618 0.0 93.646 0.163 ;
      END
   END g265666_p

   PIN g265686_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.45 0.0 94.478 0.163 ;
      END
   END g265686_p

   PIN g265687_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.194 0.0 94.222 0.163 ;
      END
   END g265687_p

   PIN g266335_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.834 0.0 86.862 0.163 ;
      END
   END g266335_p

   PIN g267264_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.554 0.0 61.582 0.163 ;
      END
   END g267264_da

   PIN g267734_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.482 0.0 66.51 0.163 ;
      END
   END g267734_p

   PIN g267768_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.33 0.0 65.358 0.163 ;
      END
   END g267768_p

   PIN g267963_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.626 0.0 64.654 0.163 ;
      END
   END g267963_p

   PIN g269325_p1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.226 0.0 106.254 0.163 ;
      END
   END g269325_p1

   PIN g270287_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.954 0.0 67.982 0.163 ;
      END
   END g270287_p

   PIN g270719_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.418 0.0 42.446 0.163 ;
      END
   END g270719_p

   PIN g270759_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.81 0.0 61.838 0.163 ;
      END
   END g270759_da

   PIN g270759_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.81 0.0 61.838 0.163 ;
      END
   END g270759_db

   PIN g271925_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.13 0.0 30.158 0.163 ;
      END
   END g271925_p

   PIN g271962_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.178 0.0 32.206 0.163 ;
      END
   END g271962_p

   PIN g271983_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.578 0.0 30.606 0.163 ;
      END
   END g271983_p

   PIN g272146_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.946 0.0 32.974 0.163 ;
      END
   END g272146_p

   PIN g273791_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.274 0.163 20.302 ;
      END
   END g273791_p

   PIN g274959_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.962 0.0 14.99 0.163 ;
      END
   END g274959_p

   PIN g275109_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.922 0.0 7.95 0.163 ;
      END
   END g275109_sb

   PIN g275315_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.202 94.557 9.23 94.72 ;
      END
   END g275315_da

   PIN g275315_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.29 94.557 10.318 94.72 ;
      END
   END g275315_db

   PIN g279718_p2
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.45 0.163 70.478 ;
      END
   END g279718_p2

   PIN g279854_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.706 0.163 62.734 ;
      END
   END g279854_p

   PIN g280604_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.994 0.163 59.022 ;
      END
   END g280604_p

   PIN g281129_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.762 0.0 3.79 0.163 ;
      END
   END g281129_p

   PIN g302688_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.778 0.0 1.806 0.163 ;
      END
   END g302688_p

   PIN g302697_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.618 0.0 5.646 0.163 ;
      END
   END g302697_p

   PIN g302698_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.698 0.163 3.726 ;
      END
   END g302698_p

   PIN g302705_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.498 0.0 8.526 0.163 ;
      END
   END g302705_p

   PIN g303296_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.442 0.163 3.47 ;
      END
   END g303296_p

   PIN g303330_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.394 0.163 9.422 ;
      END
   END g303330_p

   PIN g303332_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.49 0.0 13.518 0.163 ;
      END
   END g303332_p

   PIN g303358_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.762 0.163 3.79 ;
      END
   END g303358_p

   PIN g304265_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.802 0.0 2.83 0.163 ;
      END
   END g304265_p

   PIN g304267_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.01 0.0 9.038 0.163 ;
      END
   END g304267_p

   PIN g304295_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.21 0.0 4.238 0.163 ;
      END
   END g304295_p

   PIN g304307_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.338 0.163 20.366 ;
      END
   END g304307_p

   PIN g304312_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.226 0.0 2.254 0.163 ;
      END
   END g304312_p

   PIN g304735_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.402 0.163 12.43 ;
      END
   END g304735_p

   PIN g304777_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.458 0.163 9.486 ;
      END
   END g304777_p

   PIN g322260_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.762 0.0 67.79 0.163 ;
      END
   END g322260_p

   PIN g322487_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.45 0.0 102.478 0.163 ;
      END
   END g322487_p

   PIN g322619_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.122 0.0 51.15 0.163 ;
      END
   END g322619_da

   PIN g322619_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.378 0.0 75.406 0.163 ;
      END
   END g322619_db

   PIN n_1057
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.258 0.163 6.286 ;
      END
   END n_1057

   PIN n_108861
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.858 0.163 39.886 ;
      END
   END n_108861

   PIN n_109000
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.322 0.163 6.35 ;
      END
   END n_109000

   PIN n_109172
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.69 0.0 0.718 0.163 ;
      END
   END n_109172

   PIN n_109184
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.098 0.0 26.126 0.163 ;
      END
   END n_109184

   PIN n_1098
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.626 0.163 16.654 ;
      END
   END n_1098

   PIN n_112975
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.154 0.0 119.182 0.163 ;
      END
   END n_112975

   PIN n_112976
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.682 0.0 117.71 0.163 ;
      END
   END n_112976

   PIN n_113031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.626 0.0 72.654 0.163 ;
      END
   END n_113031

   PIN n_116915
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.842 0.0 17.87 0.163 ;
      END
   END n_116915

   PIN n_116916
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.498 0.0 8.526 0.082 ;
      END
   END n_116916

   PIN n_116953
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.69 0.0 16.718 0.163 ;
      END
   END n_116953

   PIN n_117338
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.986 0.163 8.014 ;
      END
   END n_117338

   PIN n_117342
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 5.874 0.163 5.902 ;
      END
   END n_117342

   PIN n_117601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.186 0.0 75.214 0.163 ;
      END
   END n_117601

   PIN n_117819
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.418 0.0 106.446 0.163 ;
      END
   END n_117819

   PIN n_118320
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.914 0.0 36.942 0.163 ;
      END
   END n_118320

   PIN n_118334
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.402 0.0 52.43 0.163 ;
      END
   END n_118334

   PIN n_118459
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.874 0.0 13.902 0.163 ;
      END
   END n_118459

   PIN n_118597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.682 94.557 5.71 94.72 ;
      END
   END n_118597

   PIN n_118744
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.058 0.163 59.086 ;
      END
   END n_118744

   PIN n_118754
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.698 0.0 59.726 0.163 ;
      END
   END n_118754

   PIN n_126138
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.562 0.163 16.59 ;
      END
   END n_126138

   PIN n_1264
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.29 0.0 2.318 0.163 ;
      END
   END n_1264

   PIN n_1278
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.698 0.0 3.726 0.163 ;
      END
   END n_1278

   PIN n_13895
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.298 0.0 5.326 0.163 ;
      END
   END n_13895

   PIN n_140823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.13 0.0 62.158 0.163 ;
      END
   END n_140823

   PIN n_1464
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.85 0.0 4.878 0.163 ;
      END
   END n_1464

   PIN n_1469
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.754 0.0 0.782 0.163 ;
      END
   END n_1469

   PIN n_1482
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.586 0.0 1.614 0.163 ;
      END
   END n_1482

   PIN n_1507
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 5.938 0.163 5.966 ;
      END
   END n_1507

   PIN n_1511
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.098 0.0 2.126 0.163 ;
      END
   END n_1511

   PIN n_151614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.306 0.0 0.334 0.163 ;
      END
   END n_151614

   PIN n_1599
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.082 0.163 20.11 ;
      END
   END n_1599

   PIN n_162433
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.77 0.163 62.798 ;
      END
   END n_162433

   PIN n_1790
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.466 0.163 12.494 ;
      END
   END n_1790

   PIN n_18375
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.354 0.163 66.382 ;
      END
   END n_18375

   PIN n_183956
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.61 0.0 18.638 0.163 ;
      END
   END n_183956

   PIN n_1867
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.962 0.163 6.99 ;
      END
   END n_1867

   PIN n_1932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.906 0.0 1.934 0.163 ;
      END
   END n_1932

   PIN n_1952
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.93 0.163 10.958 ;
      END
   END n_1952

   PIN n_19942
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.674 0.163 66.702 ;
      END
   END n_19942

   PIN n_19943
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.418 0.163 66.446 ;
      END
   END n_19943

   PIN n_19987
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.21 0.163 4.238 ;
      END
   END n_19987

   PIN n_20051
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.506 0.163 3.534 ;
      END
   END n_20051

   PIN n_2049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.722 0.0 4.75 0.163 ;
      END
   END n_2049

   PIN n_20823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.146 0.0 4.174 0.163 ;
      END
   END n_20823

   PIN n_20967
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.834 0.163 62.862 ;
      END
   END n_20967

   PIN n_21560
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.266 0.0 1.294 0.163 ;
      END
   END n_21560

   PIN n_21836
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.194 0.0 6.222 0.163 ;
      END
   END n_21836

   PIN n_21898
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.146 0.163 20.174 ;
      END
   END n_21898

   PIN n_21970
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.322 0.0 6.35 0.163 ;
      END
   END n_21970

   PIN n_21978
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.906 0.0 17.934 0.163 ;
      END
   END n_21978

   PIN n_21997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.818 0.0 0.846 0.163 ;
      END
   END n_21997

   PIN n_22074
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.57 0.163 11.598 ;
      END
   END n_22074

   PIN n_22077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.362 0.0 5.39 0.163 ;
      END
   END n_22077

   PIN n_22109
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.41 0.0 7.438 0.163 ;
      END
   END n_22109

   PIN n_22116
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.458 0.0 17.486 0.163 ;
      END
   END n_22116

   PIN n_22254
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.29 0.163 10.318 ;
      END
   END n_22254

   PIN n_22267
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.306 0.0 8.334 0.163 ;
      END
   END n_22267

   PIN n_22272
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.626 0.0 0.654 0.163 ;
      END
   END n_22272

   PIN n_22339
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.37 0.0 8.398 0.163 ;
      END
   END n_22339

   PIN n_22384
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.426 0.0 5.454 0.082 ;
      END
   END n_22384

   PIN n_22477
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.674 0.163 10.702 ;
      END
   END n_22477

   PIN n_22600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.522 0.0 17.55 0.163 ;
      END
   END n_22600

   PIN n_22668
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.53 0.163 12.558 ;
      END
   END n_22668

   PIN n_22760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.426 0.0 5.454 0.163 ;
      END
   END n_22760

   PIN n_22793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.554 0.0 5.582 0.163 ;
      END
   END n_22793

   PIN n_22810
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.618 0.0 5.646 0.163 ;
      END
   END n_22810

   PIN n_22832
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.434 0.163 16.462 ;
      END
   END n_22832

   PIN n_22938
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.578 0.0 6.606 0.163 ;
      END
   END n_22938

   PIN n_23072
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.042 0.0 5.07 0.163 ;
      END
   END n_23072

   PIN n_23082
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.77 0.163 6.798 ;
      END
   END n_23082

   PIN n_23089
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.034 0.163 10.062 ;
      END
   END n_23089

   PIN n_23126
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.362 0.0 5.39 0.163 ;
      END
   END n_23126

   PIN n_23209
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.146 0.0 4.174 0.163 ;
      END
   END n_23209

   PIN n_23215
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.634 0.163 11.662 ;
      END
   END n_23215

   PIN n_2327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.834 0.0 6.862 0.163 ;
      END
   END n_2327

   PIN n_23391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.066 0.0 6.094 0.163 ;
      END
   END n_23391

   PIN n_23480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.514 0.0 6.542 0.163 ;
      END
   END n_23480

   PIN n_23488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.514 0.163 6.542 ;
      END
   END n_23488

   PIN n_23559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.562 0.163 8.59 ;
      END
   END n_23559

   PIN n_23605
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.194 0.0 6.222 0.163 ;
      END
   END n_23605

   PIN n_23607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.77 0.0 6.798 0.163 ;
      END
   END n_23607

   PIN n_23658
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.346 0.0 7.374 0.163 ;
      END
   END n_23658

   PIN n_23760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.498 0.163 24.526 ;
      END
   END n_23760

   PIN n_23795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.306 0.163 8.334 ;
      END
   END n_23795

   PIN n_23805
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.21 0.163 20.238 ;
      END
   END n_23805

   PIN n_23889
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.266 94.557 129.294 94.72 ;
      END
   END n_23889

   PIN n_23929
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 167.666 0.0 167.694 0.163 ;
      END
   END n_23929

   PIN n_24160
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.738 0.163 10.766 ;
      END
   END n_24160

   PIN n_24271
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.242 0.163 24.27 ;
      END
   END n_24271

   PIN n_24308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.138 0.0 1.166 0.163 ;
      END
   END n_24308

   PIN n_24929
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.218 0.082 7.246 ;
      END
   END n_24929

   PIN n_25559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.138 0.163 9.166 ;
      END
   END n_25559

   PIN n_25809
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 81.906 0.163 81.934 ;
      END
   END n_25809

   PIN n_25811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.954 0.163 35.982 ;
      END
   END n_25811

   PIN n_25812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.898 0.163 54.926 ;
      END
   END n_25812

   PIN n_25904
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.994 0.163 3.022 ;
      END
   END n_25904

   PIN n_25932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.794 0.0 55.822 0.163 ;
      END
   END n_25932

   PIN n_25934
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 81.97 0.163 81.998 ;
      END
   END n_25934

   PIN n_25939
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.13 0.163 78.158 ;
      END
   END n_25939

   PIN n_25994
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.562 0.163 24.59 ;
      END
   END n_25994

   PIN n_26053
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 89.522 0.163 89.55 ;
      END
   END n_26053

   PIN n_26162
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.018 0.0 4.046 0.163 ;
      END
   END n_26162

   PIN n_26171
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.962 0.082 14.99 ;
      END
   END n_26171

   PIN n_26172
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.938 0.163 13.966 ;
      END
   END n_26172

   PIN n_26188
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.034 0.163 82.062 ;
      END
   END n_26188

   PIN n_26255
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.258 0.163 14.286 ;
      END
   END n_26255

   PIN n_26333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.418 0.0 2.446 0.163 ;
      END
   END n_26333

   PIN n_26360
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.93 0.163 2.958 ;
      END
   END n_26360

   PIN n_26362
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.402 0.163 20.43 ;
      END
   END n_26362

   PIN n_26373
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.09 0.163 15.118 ;
      END
   END n_26373

   PIN n_26495
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.45 0.163 14.478 ;
      END
   END n_26495

   PIN n_26507
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.122 0.163 3.15 ;
      END
   END n_26507

   PIN n_26533
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.066 0.163 14.094 ;
      END
   END n_26533

   PIN n_26619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.114 0.163 8.142 ;
      END
   END n_26619

   PIN n_26627
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.986 0.163 16.014 ;
      END
   END n_26627

   PIN n_26634
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.986 0.163 32.014 ;
      END
   END n_26634

   PIN n_26662
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.154 0.163 15.182 ;
      END
   END n_26662

   PIN n_26750
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.466 0.163 20.494 ;
      END
   END n_26750

   PIN n_26760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.514 0.163 14.542 ;
      END
   END n_26760

   PIN n_26773
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.018 0.163 20.046 ;
      END
   END n_26773

   PIN n_26775
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 13.234 0.163 13.262 ;
      END
   END n_26775

   PIN n_26929
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.898 0.163 6.926 ;
      END
   END n_26929

   PIN n_27125
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.946 0.0 24.974 0.163 ;
      END
   END n_27125

   PIN n_27252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.178 0.163 8.206 ;
      END
   END n_27252

   PIN n_27259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.578 0.163 14.606 ;
      END
   END n_27259

   PIN n_27388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.762 0.163 11.79 ;
      END
   END n_27388

   PIN n_27391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.378 0.163 3.406 ;
      END
   END n_27391

   PIN n_27437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.41 0.163 15.438 ;
      END
   END n_27437

   PIN n_27439
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.49 0.0 29.518 0.163 ;
      END
   END n_27439

   PIN n_27513
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.746 94.557 21.774 94.72 ;
      END
   END n_27513

   PIN n_2774
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.954 0.0 3.982 0.163 ;
      END
   END n_2774

   PIN n_27816
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.418 0.0 34.446 0.163 ;
      END
   END n_27816

   PIN n_27849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.386 0.0 6.414 0.163 ;
      END
   END n_27849

   PIN n_27887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.794 0.0 55.822 0.163 ;
      END
   END n_27887

   PIN n_27899
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.754 0.0 24.782 0.163 ;
      END
   END n_27899

   PIN n_27900
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.818 0.0 48.846 0.163 ;
      END
   END n_27900

   PIN n_27929
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.266 0.0 33.294 0.163 ;
      END
   END n_27929

   PIN n_27947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.298 0.0 13.326 0.163 ;
      END
   END n_27947

   PIN n_27948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.33 0.0 33.358 0.163 ;
      END
   END n_27948

   PIN n_28029
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.626 0.0 32.654 0.163 ;
      END
   END n_28029

   PIN n_28094
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.634 0.0 59.662 0.163 ;
      END
   END n_28094

   PIN n_28111
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.65 0.0 33.678 0.163 ;
      END
   END n_28111

   PIN n_28189
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.538 0.0 31.566 0.163 ;
      END
   END n_28189

   PIN n_28201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.434 0.0 32.462 0.163 ;
      END
   END n_28201

   PIN n_28213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.946 0.0 40.974 0.163 ;
      END
   END n_28213

   PIN n_28224
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.106 0.0 61.134 0.163 ;
      END
   END n_28224

   PIN n_28276
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.066 0.0 62.094 0.163 ;
      END
   END n_28276

   PIN n_28296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.57 0.0 59.598 0.163 ;
      END
   END n_28296

   PIN n_28297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.914 0.0 60.942 0.163 ;
      END
   END n_28297

   PIN n_28299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.754 0.0 64.782 0.163 ;
      END
   END n_28299

   PIN n_28326
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.786 0.0 20.814 0.163 ;
      END
   END n_28326

   PIN n_28348
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.394 0.0 33.422 0.163 ;
      END
   END n_28348

   PIN n_28350
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.658 0.0 36.686 0.163 ;
      END
   END n_28350

   PIN n_28372
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.25 0.0 59.278 0.163 ;
      END
   END n_28372

   PIN n_28387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.17 0.0 37.198 0.163 ;
      END
   END n_28387

   PIN n_28388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.234 0.0 37.262 0.163 ;
      END
   END n_28388

   PIN n_28399
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.01 0.0 65.038 0.163 ;
      END
   END n_28399

   PIN n_28430
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.434 0.0 32.462 0.163 ;
      END
   END n_28430

   PIN n_28431
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.874 0.0 29.902 0.163 ;
      END
   END n_28431

   PIN n_28457
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.93 0.0 58.958 0.163 ;
      END
   END n_28457

   PIN n_28473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.818 0.0 64.846 0.163 ;
      END
   END n_28473

   PIN n_28474
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.818 0.0 56.846 0.163 ;
      END
   END n_28474

   PIN n_28500
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.266 0.0 65.294 0.163 ;
      END
   END n_28500

   PIN n_28511
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.938 0.0 29.966 0.163 ;
      END
   END n_28511

   PIN n_28582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.122 0.0 59.15 0.163 ;
      END
   END n_28582

   PIN n_28583
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.682 0.0 61.71 0.163 ;
      END
   END n_28583

   PIN n_28596
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.226 0.0 66.254 0.163 ;
      END
   END n_28596

   PIN n_28623
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.074 0.0 33.102 0.163 ;
      END
   END n_28623

   PIN n_28722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.554 0.0 29.582 0.163 ;
      END
   END n_28722

   PIN n_28734
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.906 0.0 65.934 0.163 ;
      END
   END n_28734

   PIN n_28743
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.69 0.0 64.718 0.163 ;
      END
   END n_28743

   PIN n_28749
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.714 0.0 25.742 0.163 ;
      END
   END n_28749

   PIN n_28755
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.066 0.0 62.094 0.163 ;
      END
   END n_28755

   PIN n_28760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.89 0.0 59.918 0.163 ;
      END
   END n_28760

   PIN n_28763
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.994 0.0 59.022 0.163 ;
      END
   END n_28763

   PIN n_28782
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.298 0.0 37.326 0.163 ;
      END
   END n_28782

   PIN n_28794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.706 0.0 6.734 0.163 ;
      END
   END n_28794

   PIN n_28827
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.074 0.0 41.102 0.163 ;
      END
   END n_28827

   PIN n_28860
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.466 0.0 60.494 0.163 ;
      END
   END n_28860

   PIN n_28864
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.714 0.0 33.742 0.163 ;
      END
   END n_28864

   PIN n_28869
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.306 0.0 32.334 0.163 ;
      END
   END n_28869

   PIN n_28888
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.458 0.0 33.486 0.163 ;
      END
   END n_28888

   PIN n_28929
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.73 0.0 31.758 0.163 ;
      END
   END n_28929

   PIN n_28938
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.938 0.0 29.966 0.163 ;
      END
   END n_28938

   PIN n_28986
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.978 0.0 37.006 0.163 ;
      END
   END n_28986

   PIN n_29006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.242 0.0 32.27 0.163 ;
      END
   END n_29006

   PIN n_29039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.85 0.0 36.878 0.163 ;
      END
   END n_29039

   PIN n_29060
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.594 0.0 36.622 0.163 ;
      END
   END n_29060

   PIN n_29083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.818 0.0 32.846 0.163 ;
      END
   END n_29083

   PIN n_29086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.962 0.0 30.99 0.163 ;
      END
   END n_29086

   PIN n_29128
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.154 0.0 31.182 0.163 ;
      END
   END n_29128

   PIN n_29133
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.418 0.0 58.446 0.163 ;
      END
   END n_29133

   PIN n_29140
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.802 0.0 58.83 0.163 ;
      END
   END n_29140

   PIN n_29154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.042 0.0 37.07 0.163 ;
      END
   END n_29154

   PIN n_29251
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.498 0.0 32.526 0.163 ;
      END
   END n_29251

   PIN n_29269
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.41 0.0 31.438 0.163 ;
      END
   END n_29269

   PIN n_29329
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.354 0.0 42.382 0.163 ;
      END
   END n_29329

   PIN n_29418
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.362 0.0 37.39 0.163 ;
      END
   END n_29418

   PIN n_29426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.426 0.0 37.454 0.163 ;
      END
   END n_29426

   PIN n_29527
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 57.202 0.0 57.23 0.163 ;
      END
   END n_29527

   PIN n_29608
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.434 0.0 56.462 0.163 ;
      END
   END n_29608

   PIN n_29625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.106 0.0 37.134 0.163 ;
      END
   END n_29625

   PIN n_29647
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.578 0.0 54.606 0.163 ;
      END
   END n_29647

   PIN n_29648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.682 0.0 29.71 0.163 ;
      END
   END n_29648

   PIN n_29650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.874 0.0 29.902 0.163 ;
      END
   END n_29650

   PIN n_29674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.298 0.0 29.326 0.163 ;
      END
   END n_29674

   PIN n_29692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.33 0.0 121.358 0.163 ;
      END
   END n_29692

   PIN n_29701
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.962 0.0 54.99 0.163 ;
      END
   END n_29701

   PIN n_29719
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.522 0.0 33.55 0.163 ;
      END
   END n_29719

   PIN n_29721
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.514 0.0 102.542 0.163 ;
      END
   END n_29721

   PIN n_29723
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.218 0.0 55.246 0.163 ;
      END
   END n_29723

   PIN n_29738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.178 0.0 56.206 0.163 ;
      END
   END n_29738

   PIN n_29760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.778 0.0 113.806 0.163 ;
      END
   END n_29760

   PIN n_29815
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.082 0.0 52.11 0.163 ;
      END
   END n_29815

   PIN n_29847
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.666 0.0 31.694 0.163 ;
      END
   END n_29847

   PIN n_29871
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.002 0.0 54.03 0.163 ;
      END
   END n_29871

   PIN n_29888
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.49 0.0 61.518 0.163 ;
      END
   END n_29888

   PIN n_2989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.498 0.163 16.526 ;
      END
   END n_2989

   PIN n_30044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.866 0.0 106.894 0.163 ;
      END
   END n_30044

   PIN n_3007
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.754 0.163 8.782 ;
      END
   END n_3007

   PIN n_30077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.514 0.0 118.542 0.163 ;
      END
   END n_30077

   PIN n_30138
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.41 0.0 71.438 0.163 ;
      END
   END n_30138

   PIN n_30169
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.666 0.0 119.694 0.163 ;
      END
   END n_30169

   PIN n_30172
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.442 0.0 107.47 0.163 ;
      END
   END n_30172

   PIN n_30223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.522 0.0 113.55 0.163 ;
      END
   END n_30223

   PIN n_30282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.09 0.0 119.118 0.163 ;
      END
   END n_30282

   PIN n_30287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.114 0.0 104.142 0.163 ;
      END
   END n_30287

   PIN n_30333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.53 0.0 36.558 0.163 ;
      END
   END n_30333

   PIN n_30356
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.362 0.0 109.39 0.163 ;
      END
   END n_30356

   PIN n_30360
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.202 0.0 129.23 0.163 ;
      END
   END n_30360

   PIN n_30370
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.946 0.0 136.974 0.163 ;
      END
   END n_30370

   PIN n_30373
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.522 0.0 121.55 0.163 ;
      END
   END n_30373

   PIN n_30387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.986 0.0 120.014 0.163 ;
      END
   END n_30387

   PIN n_30388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.794 0.0 119.822 0.163 ;
      END
   END n_30388

   PIN n_30391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.722 0.0 116.75 0.163 ;
      END
   END n_30391

   PIN n_30392
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.146 0.0 116.174 0.163 ;
      END
   END n_30392

   PIN n_30407
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.954 0.0 107.982 0.163 ;
      END
   END n_30407

   PIN n_30426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.17 0.0 117.198 0.163 ;
      END
   END n_30426

   PIN n_30437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.362 0.0 125.39 0.163 ;
      END
   END n_30437

   PIN n_30480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.602 0.0 119.63 0.163 ;
      END
   END n_30480

   PIN n_30487
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.954 0.0 35.982 0.163 ;
      END
   END n_30487

   PIN n_30496
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.754 0.0 40.782 0.163 ;
      END
   END n_30496

   PIN n_30609
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.082 0.0 116.11 0.163 ;
      END
   END n_30609

   PIN n_30616
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 68.018 0.0 68.046 0.163 ;
      END
   END n_30616

   PIN n_30646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.05 0.0 104.078 0.163 ;
      END
   END n_30646

   PIN n_30656
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.49 0.0 109.518 0.163 ;
      END
   END n_30656

   PIN n_30667
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.762 0.0 115.79 0.163 ;
      END
   END n_30667

   PIN n_30673
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.426 0.0 117.454 0.163 ;
      END
   END n_30673

   PIN n_30685
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 133.042 0.0 133.07 0.163 ;
      END
   END n_30685

   PIN n_30712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.61 0.0 106.638 0.163 ;
      END
   END n_30712

   PIN n_30782
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.618 0.0 109.646 0.163 ;
      END
   END n_30782

   PIN n_30795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.81 0.0 109.838 0.163 ;
      END
   END n_30795

   PIN n_30846
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.658 0.0 116.686 0.163 ;
      END
   END n_30846

   PIN n_30872
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.914 0.0 116.942 0.163 ;
      END
   END n_30872

   PIN n_30945
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.602 0.0 63.63 0.163 ;
      END
   END n_30945

   PIN n_30958
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.906 0.0 113.934 0.163 ;
      END
   END n_30958

   PIN n_30959
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.146 0.0 108.174 0.163 ;
      END
   END n_30959

   PIN n_30977
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.89 0.0 67.918 0.163 ;
      END
   END n_30977

   PIN n_30991
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.098 0.0 106.126 0.163 ;
      END
   END n_30991

   PIN n_31042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.554 0.0 117.582 0.163 ;
      END
   END n_31042

   PIN n_31076
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.874 0.0 109.902 0.163 ;
      END
   END n_31076

   PIN n_31092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.706 0.0 110.734 0.163 ;
      END
   END n_31092

   PIN n_31119
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.778 0.0 105.806 0.163 ;
      END
   END n_31119

   PIN n_31120
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.554 0.0 109.582 0.082 ;
      END
   END n_31120

   PIN n_31170
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.258 0.0 110.286 0.163 ;
      END
   END n_31170

   PIN n_31173
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.842 0.0 105.87 0.163 ;
      END
   END n_31173

   PIN n_31184
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.746 0.0 109.774 0.163 ;
      END
   END n_31184

   PIN n_31185
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.682 0.0 109.71 0.163 ;
      END
   END n_31185

   PIN n_31195
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.874 0.0 109.902 0.163 ;
      END
   END n_31195

   PIN n_31218
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.938 0.0 109.966 0.163 ;
      END
   END n_31218

   PIN n_31239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.186 0.0 115.214 0.163 ;
      END
   END n_31239

   PIN n_31271
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.322 0.0 110.35 0.163 ;
      END
   END n_31271

   PIN n_31355
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.906 0.0 105.934 0.163 ;
      END
   END n_31355

   PIN n_31403
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.786 0.0 108.814 0.163 ;
      END
   END n_31403

   PIN n_31424
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.882 0.0 104.91 0.163 ;
      END
   END n_31424

   PIN n_31460
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.298 0.0 109.326 0.163 ;
      END
   END n_31460

   PIN n_31476
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.57 0.0 115.598 0.163 ;
      END
   END n_31476

   PIN n_31484
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.498 0.0 40.526 0.163 ;
      END
   END n_31484

   PIN n_31490
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.722 0.0 108.75 0.163 ;
      END
   END n_31490

   PIN n_31494
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.786 0.0 108.814 0.163 ;
      END
   END n_31494

   PIN n_31516
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.29 0.0 114.318 0.163 ;
      END
   END n_31516

   PIN n_3166
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.826 0.163 3.854 ;
      END
   END n_3166

   PIN n_31689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.306 0.0 112.334 0.163 ;
      END
   END n_31689

   PIN n_31709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.218 0.0 111.246 0.163 ;
      END
   END n_31709

   PIN n_31727
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.042 0.0 101.07 0.163 ;
      END
   END n_31727

   PIN n_31730
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.786 0.0 44.814 0.163 ;
      END
   END n_31730

   PIN n_31731
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.122 0.0 19.15 0.163 ;
      END
   END n_31731

   PIN n_31732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.706 0.0 110.734 0.163 ;
      END
   END n_31732

   PIN n_31734
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.666 0.0 47.694 0.163 ;
      END
   END n_31734

   PIN n_31751
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.354 0.0 98.382 0.163 ;
      END
   END n_31751

   PIN n_31856
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.25 0.0 75.278 0.163 ;
      END
   END n_31856

   PIN n_31919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.714 0.0 73.742 0.163 ;
      END
   END n_31919

   PIN n_32004
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.834 0.0 70.862 0.163 ;
      END
   END n_32004

   PIN n_32213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.234 0.0 69.262 0.163 ;
      END
   END n_32213

   PIN n_32267
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.21 0.0 68.238 0.163 ;
      END
   END n_32267

   PIN n_32307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.602 0.0 71.63 0.163 ;
      END
   END n_32307

   PIN n_32336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.53 0.0 68.558 0.163 ;
      END
   END n_32336

   PIN n_32337
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.57 0.0 75.598 0.163 ;
      END
   END n_32337

   PIN n_32344
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.506 0.0 67.534 0.163 ;
      END
   END n_32344

   PIN n_32386
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.706 0.0 70.734 0.163 ;
      END
   END n_32386

   PIN n_32387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.938 0.0 69.966 0.163 ;
      END
   END n_32387

   PIN n_32400
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.778 0.0 41.806 0.163 ;
      END
   END n_32400

   PIN n_32435
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.858 0.0 71.886 0.163 ;
      END
   END n_32435

   PIN n_32665
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.402 0.0 52.43 0.163 ;
      END
   END n_32665

   PIN n_32697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.466 0.0 52.494 0.163 ;
      END
   END n_32697

   PIN n_32701
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.722 0.0 68.75 0.163 ;
      END
   END n_32701

   PIN n_32779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.634 0.0 67.662 0.163 ;
      END
   END n_32779

   PIN n_32785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.826 0.0 67.854 0.163 ;
      END
   END n_32785

   PIN n_32805
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.41 0.0 71.438 0.163 ;
      END
   END n_32805

   PIN n_32833
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.634 0.0 75.662 0.163 ;
      END
   END n_32833

   PIN n_32842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.474 0.0 71.502 0.163 ;
      END
   END n_32842

   PIN n_32845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.442 0.0 75.47 0.163 ;
      END
   END n_32845

   PIN n_32893
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.026 0.0 71.054 0.163 ;
      END
   END n_32893

   PIN n_32923
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.498 0.0 48.526 0.163 ;
      END
   END n_32923

   PIN n_32979
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.778 0.0 65.806 0.163 ;
      END
   END n_32979

   PIN n_3304
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.098 0.0 2.126 0.163 ;
      END
   END n_3304

   PIN n_33066
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.082 0.0 52.11 0.163 ;
      END
   END n_33066

   PIN n_33072
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.41 0.0 63.438 0.163 ;
      END
   END n_33072

   PIN n_33082
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.314 0.0 75.342 0.163 ;
      END
   END n_33082

   PIN n_33099
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.826 0.0 67.854 0.163 ;
      END
   END n_33099

   PIN n_33111
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.858 0.0 55.886 0.163 ;
      END
   END n_33111

   PIN n_33201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.858 0.0 55.886 0.163 ;
      END
   END n_33201

   PIN n_33206
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.762 0.0 59.79 0.163 ;
      END
   END n_33206

   PIN n_33211
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.474 0.0 63.502 0.163 ;
      END
   END n_33211

   PIN n_33227
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.602 0.0 63.63 0.163 ;
      END
   END n_33227

   PIN n_33245
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.546 0.0 66.574 0.163 ;
      END
   END n_33245

   PIN n_33253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 72.114 0.0 72.142 0.163 ;
      END
   END n_33253

   PIN n_33287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.314 0.0 59.342 0.163 ;
      END
   END n_33287

   PIN n_33296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 68.146 0.0 68.174 0.163 ;
      END
   END n_33296

   PIN n_33327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.642 0.0 70.67 0.163 ;
      END
   END n_33327

   PIN n_33328
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.666 0.0 63.694 0.163 ;
      END
   END n_33328

   PIN n_33329
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.73 0.0 63.758 0.163 ;
      END
   END n_33329

   PIN n_33422
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.37 0.0 48.398 0.163 ;
      END
   END n_33422

   PIN n_33463
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.922 0.0 55.95 0.163 ;
      END
   END n_33463

   PIN n_33484
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 80.69 0.0 80.718 0.163 ;
      END
   END n_33484

   PIN n_3349
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.386 0.163 6.414 ;
      END
   END n_3349

   PIN n_33490
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.562 0.0 48.59 0.163 ;
      END
   END n_33490

   PIN n_33562
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.45 0.0 62.478 0.163 ;
      END
   END n_33562

   PIN n_33566
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.034 0.0 66.062 0.163 ;
      END
   END n_33566

   PIN n_33587
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.538 0.0 63.566 0.163 ;
      END
   END n_33587

   PIN n_33588
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.498 0.0 64.526 0.163 ;
      END
   END n_33588

   PIN n_33614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.61 0.0 42.638 0.163 ;
      END
   END n_33614

   PIN n_33630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.146 0.0 52.174 0.163 ;
      END
   END n_33630

   PIN n_3365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.594 0.163 12.622 ;
      END
   END n_3365

   PIN n_33653
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.986 0.0 56.014 0.163 ;
      END
   END n_33653

   PIN n_33655
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.922 0.0 55.95 0.163 ;
      END
   END n_33655

   PIN n_33657
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.21 0.0 52.238 0.163 ;
      END
   END n_33657

   PIN n_33686
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.626 94.557 144.654 94.72 ;
      END
   END n_33686

   PIN n_33750
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 133.106 0.0 133.134 0.163 ;
      END
   END n_33750

   PIN n_33757
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.122 0.0 83.15 0.163 ;
      END
   END n_33757

   PIN n_34020
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.738 0.0 90.766 0.163 ;
      END
   END n_34020

   PIN n_34137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.09 0.0 87.118 0.163 ;
      END
   END n_34137

   PIN n_34143
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.57 0.0 91.598 0.163 ;
      END
   END n_34143

   PIN n_34216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.314 0.0 91.342 0.163 ;
      END
   END n_34216

   PIN n_34299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.154 0.0 87.182 0.163 ;
      END
   END n_34299

   PIN n_34438
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.426 0.0 93.454 0.163 ;
      END
   END n_34438

   PIN n_34477
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.738 0.0 90.766 0.082 ;
      END
   END n_34477

   PIN n_34478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.73 0.0 63.758 0.163 ;
      END
   END n_34478

   PIN n_34489
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.122 0.0 91.15 0.163 ;
      END
   END n_34489

   PIN n_34500
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.186 0.0 91.214 0.163 ;
      END
   END n_34500

   PIN n_34748
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.346 0.0 95.374 0.163 ;
      END
   END n_34748

   PIN n_34749
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.962 0.0 94.99 0.163 ;
      END
   END n_34749

   PIN n_34758
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.906 0.0 89.934 0.163 ;
      END
   END n_34758

   PIN n_34759
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.61 0.0 90.638 0.163 ;
      END
   END n_34759

   PIN n_34760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.21 0.0 92.238 0.163 ;
      END
   END n_34760

   PIN n_34775
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.634 0.0 91.662 0.163 ;
      END
   END n_34775

   PIN n_34788
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.898 0.0 86.926 0.163 ;
      END
   END n_34788

   PIN n_3487
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.002 0.163 6.03 ;
      END
   END n_3487

   PIN n_34902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.018 0.0 92.046 0.163 ;
      END
   END n_34902

   PIN n_34904
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.514 0.0 94.542 0.163 ;
      END
   END n_34904

   PIN n_34943
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.298 0.0 93.326 0.163 ;
      END
   END n_34943

   PIN n_35025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.322 0.0 94.35 0.163 ;
      END
   END n_35025

   PIN n_35036
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.682 0.0 93.71 0.163 ;
      END
   END n_35036

   PIN n_35105
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.258 0.0 94.286 0.163 ;
      END
   END n_35105

   PIN n_35129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.25 0.0 91.278 0.163 ;
      END
   END n_35129

   PIN n_35131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.714 0.0 89.742 0.163 ;
      END
   END n_35131

   PIN n_35134
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.554 0.0 93.582 0.163 ;
      END
   END n_35134

   PIN n_35140
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.61 0.0 90.638 0.163 ;
      END
   END n_35140

   PIN n_35143
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.698 0.0 91.726 0.163 ;
      END
   END n_35143

   PIN n_35375
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 87.09 0.0 87.118 0.163 ;
      END
   END n_35375

   PIN n_35580
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.77 0.0 94.798 0.163 ;
      END
   END n_35580

   PIN n_4090
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.354 0.163 10.382 ;
      END
   END n_4090

   PIN n_4133
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.578 0.0 6.606 0.163 ;
      END
   END n_4133

   PIN n_4333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.33 0.0 1.358 0.163 ;
      END
   END n_4333

   PIN n_4413
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.61 0.0 10.638 0.163 ;
      END
   END n_4413

   PIN n_4526
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.066 0.163 6.094 ;
      END
   END n_4526

   PIN n_4634
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.194 0.163 78.222 ;
      END
   END n_4634

   PIN n_4673
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.05 0.163 32.078 ;
      END
   END n_4673

   PIN n_4761
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.89 0.163 3.918 ;
      END
   END n_4761

   PIN n_4889
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.13 0.163 6.158 ;
      END
   END n_4889

   PIN n_4902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 85.682 0.163 85.71 ;
      END
   END n_4902

   PIN n_4922
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.53 0.163 20.558 ;
      END
   END n_4922

   PIN n_5077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.45 0.163 6.478 ;
      END
   END n_5077

   PIN n_62095
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.37 0.163 8.398 ;
      END
   END n_62095

   PIN n_63235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.522 0.163 9.55 ;
      END
   END n_63235

   PIN n_63270
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.418 0.163 10.446 ;
      END
   END n_63270

   PIN n_63281
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.962 0.0 6.99 0.163 ;
      END
   END n_63281

   PIN n_63816
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.754 0.0 24.782 0.163 ;
      END
   END n_63816

   PIN n_64050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.666 0.0 23.694 0.163 ;
      END
   END n_64050

   PIN n_64089
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.37 0.0 24.398 0.163 ;
      END
   END n_64089

   PIN n_64141
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.114 0.0 24.142 0.163 ;
      END
   END n_64141

   PIN n_64164
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.778 0.0 25.806 0.163 ;
      END
   END n_64164

   PIN n_64228
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.282 0.0 23.31 0.163 ;
      END
   END n_64228

   PIN n_64301
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.106 0.0 21.134 0.163 ;
      END
   END n_64301

   PIN n_64325
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.402 0.0 20.43 0.163 ;
      END
   END n_64325

   PIN n_64384
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.922 0.0 23.95 0.163 ;
      END
   END n_64384

   PIN n_64437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.73 0.0 23.758 0.163 ;
      END
   END n_64437

   PIN n_64570
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.002 0.0 22.03 0.163 ;
      END
   END n_64570

   PIN n_64704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.842 0.0 25.87 0.163 ;
      END
   END n_64704

   PIN n_64735
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.474 0.0 23.502 0.163 ;
      END
   END n_64735

   PIN n_64770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.57 0.163 43.598 ;
      END
   END n_64770

   PIN n_64800
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.618 0.0 21.646 0.163 ;
      END
   END n_64800

   PIN n_64801
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.21 0.0 20.238 0.163 ;
      END
   END n_64801

   PIN n_64811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.898 0.163 62.926 ;
      END
   END n_64811

   PIN n_64946
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.826 0.0 19.854 0.163 ;
      END
   END n_64946

   PIN n_64982
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.25 0.0 19.278 0.163 ;
      END
   END n_64982

   PIN n_65063
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.314 0.0 19.342 0.163 ;
      END
   END n_65063

   PIN n_65156
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.594 0.0 20.622 0.163 ;
      END
   END n_65156

   PIN n_65198
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.338 0.0 20.366 0.163 ;
      END
   END n_65198

   PIN n_65585
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.186 0.0 27.214 0.163 ;
      END
   END n_65585

   PIN n_65644
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.698 0.163 3.726 ;
      END
   END n_65644

   PIN n_65659
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.402 94.557 52.43 94.72 ;
      END
   END n_65659

   PIN n_65667
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.97 0.0 25.998 0.163 ;
      END
   END n_65667

   PIN n_65746
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.762 0.163 3.79 ;
      END
   END n_65746

   PIN n_65780
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.026 0.0 15.054 0.163 ;
      END
   END n_65780

   PIN n_65811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.186 0.163 3.214 ;
      END
   END n_65811

   PIN n_65824
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.626 0.0 16.654 0.163 ;
      END
   END n_65824

   PIN n_65827
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.466 94.557 52.494 94.72 ;
      END
   END n_65827

   PIN n_65830
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.594 0.163 12.622 ;
      END
   END n_65830

   PIN n_65889
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.41 0.163 39.438 ;
      END
   END n_65889

   PIN n_65900
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.89 0.0 27.918 0.163 ;
      END
   END n_65900

   PIN n_65921
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.738 0.0 26.766 0.163 ;
      END
   END n_65921

   PIN n_65938
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.154 0.0 15.182 0.163 ;
      END
   END n_65938

   PIN n_65939
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.322 0.0 14.35 0.163 ;
      END
   END n_65939

   PIN n_65940
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.354 0.163 10.382 ;
      END
   END n_65940

   PIN n_65963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.018 0.0 28.046 0.163 ;
      END
   END n_65963

   PIN n_66043
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.77 0.0 14.798 0.163 ;
      END
   END n_66043

   PIN n_66049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.258 0.0 14.286 0.163 ;
      END
   END n_66049

   PIN n_66062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.402 0.163 12.43 ;
      END
   END n_66062

   PIN n_66063
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.018 0.163 36.046 ;
      END
   END n_66063

   PIN n_66064
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.634 0.163 35.662 ;
      END
   END n_66064

   PIN n_66072
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.698 0.0 27.726 0.163 ;
      END
   END n_66072

   PIN n_66147
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.762 0.0 11.79 0.163 ;
      END
   END n_66147

   PIN n_66148
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.834 0.0 14.862 0.163 ;
      END
   END n_66148

   PIN n_66150
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.418 0.0 26.446 0.163 ;
      END
   END n_66150

   PIN n_66151
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.618 0.0 29.646 0.163 ;
      END
   END n_66151

   PIN n_66163
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.202 0.163 9.23 ;
      END
   END n_66163

   PIN n_66220
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.33 0.0 25.358 0.163 ;
      END
   END n_66220

   PIN n_66234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.226 0.163 10.254 ;
      END
   END n_66234

   PIN n_66256
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.506 0.0 27.534 0.163 ;
      END
   END n_66256

   PIN n_66277
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.658 0.163 12.686 ;
      END
   END n_66277

   PIN n_66320
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.586 94.557 25.614 94.72 ;
      END
   END n_66320

   PIN n_66322
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.122 0.0 27.15 0.163 ;
      END
   END n_66322

   PIN n_66366
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.57 0.163 35.598 ;
      END
   END n_66366

   PIN n_66379
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.826 0.163 3.854 ;
      END
   END n_66379

   PIN n_66409
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.21 0.0 28.238 0.163 ;
      END
   END n_66409

   PIN n_66421
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.722 0.163 12.75 ;
      END
   END n_66421

   PIN n_66434
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.786 0.163 12.814 ;
      END
   END n_66434

   PIN n_66456
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.138 0.0 25.166 0.163 ;
      END
   END n_66456

   PIN n_66462
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.346 0.163 7.374 ;
      END
   END n_66462

   PIN n_66488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.018 0.163 12.046 ;
      END
   END n_66488

   PIN n_66520
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.282 0.0 7.31 0.082 ;
      END
   END n_66520

   PIN n_66544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.042 0.0 13.07 0.163 ;
      END
   END n_66544

   PIN n_66548
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.586 0.0 25.614 0.163 ;
      END
   END n_66548

   PIN n_66565
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.962 0.0 6.99 0.163 ;
      END
   END n_66565

   PIN n_66570
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.818 0.163 8.846 ;
      END
   END n_66570

   PIN n_66577
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.21 0.163 12.238 ;
      END
   END n_66577

   PIN n_66582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.018 0.0 28.046 0.163 ;
      END
   END n_66582

   PIN n_66586
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.026 0.0 7.054 0.163 ;
      END
   END n_66586

   PIN n_66593
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.162 0.0 26.19 0.163 ;
      END
   END n_66593

   PIN n_66595
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.13 0.0 14.158 0.163 ;
      END
   END n_66595

   PIN n_66622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.85 0.163 12.878 ;
      END
   END n_66622

   PIN n_66638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.09 0.0 7.118 0.163 ;
      END
   END n_66638

   PIN n_66647
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.45 0.0 14.478 0.163 ;
      END
   END n_66647

   PIN n_66650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.802 0.0 26.83 0.163 ;
      END
   END n_66650

   PIN n_66655
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.082 0.163 36.11 ;
      END
   END n_66655

   PIN n_66706
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.194 0.163 6.222 ;
      END
   END n_66706

   PIN n_66765
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.658 0.163 12.686 ;
      END
   END n_66765

   PIN n_66766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.994 0.163 11.022 ;
      END
   END n_66766

   PIN n_66777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.186 0.0 27.214 0.163 ;
      END
   END n_66777

   PIN n_66845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.338 0.0 12.366 0.163 ;
      END
   END n_66845

   PIN n_66858
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.65 0.0 25.678 0.163 ;
      END
   END n_66858

   PIN n_66866
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.442 0.163 43.47 ;
      END
   END n_66866

   PIN n_66877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.082 0.163 12.11 ;
      END
   END n_66877

   PIN n_66939
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.506 0.163 43.534 ;
      END
   END n_66939

   PIN n_66996
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.17 0.0 21.198 0.163 ;
      END
   END n_66996

   PIN n_67014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.226 0.0 26.254 0.163 ;
      END
   END n_67014

   PIN n_67059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.106 0.0 13.134 0.163 ;
      END
   END n_67059

   PIN n_67072
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.57 0.0 11.598 0.163 ;
      END
   END n_67072

   PIN n_67086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.722 0.163 12.75 ;
      END
   END n_67086

   PIN n_67110
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.474 0.163 39.502 ;
      END
   END n_67110

   PIN n_67204
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.21 0.0 4.238 0.163 ;
      END
   END n_67204

   PIN n_67239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.378 0.0 3.406 0.163 ;
      END
   END n_67239

   PIN n_67252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.178 0.0 0.206 0.163 ;
      END
   END n_67252

   PIN n_67253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.314 0.0 11.342 0.163 ;
      END
   END n_67253

   PIN n_67287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.594 0.163 20.622 ;
      END
   END n_67287

   PIN n_6732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.554 0.0 53.582 0.163 ;
      END
   END n_6732

   PIN n_67320
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.618 0.0 13.646 0.163 ;
      END
   END n_67320

   PIN n_67524
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.706 0.0 14.734 0.163 ;
      END
   END n_67524

   PIN n_67561
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.226 0.0 18.254 0.163 ;
      END
   END n_67561

   PIN n_67606
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.682 0.0 29.71 0.163 ;
      END
   END n_67606

   PIN n_67801
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.714 0.0 17.742 0.163 ;
      END
   END n_67801

   PIN n_67898
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.906 0.0 25.934 0.163 ;
      END
   END n_67898

   PIN n_67995
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.354 0.0 18.382 0.163 ;
      END
   END n_67995

   PIN n_68021
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.266 0.0 17.294 0.163 ;
      END
   END n_68021

   PIN n_68043
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.946 0.0 16.974 0.163 ;
      END
   END n_68043

   PIN n_68092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.242 0.0 16.27 0.163 ;
      END
   END n_68092

   PIN n_68186
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.778 0.0 17.806 0.163 ;
      END
   END n_68186

   PIN n_68213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.042 0.0 21.07 0.163 ;
      END
   END n_68213

   PIN n_68361
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.034 0.0 18.062 0.163 ;
      END
   END n_68361

   PIN n_68364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.058 0.0 19.086 0.163 ;
      END
   END n_68364

   PIN n_68492
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.394 0.0 17.422 0.163 ;
      END
   END n_68492

   PIN n_68493
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.202 0.0 17.23 0.163 ;
      END
   END n_68493

   PIN n_68509
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.138 0.0 17.166 0.163 ;
      END
   END n_68509

   PIN n_68549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.418 0.0 18.446 0.163 ;
      END
   END n_68549

   PIN n_68730
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.002 0.0 30.03 0.163 ;
      END
   END n_68730

   PIN n_68839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.01 0.0 17.038 0.163 ;
      END
   END n_68839

   PIN n_68842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.074 0.0 17.102 0.163 ;
      END
   END n_68842

   PIN n_69233
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.594 0.0 12.622 0.163 ;
      END
   END n_69233

   PIN n_69250
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.73 0.0 7.758 0.163 ;
      END
   END n_69250

   PIN n_69476
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.426 0.0 109.454 0.163 ;
      END
   END n_69476

   PIN n_69494
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.722 0.0 20.75 0.163 ;
      END
   END n_69494

   PIN n_69523
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.354 0.0 98.382 0.163 ;
      END
   END n_69523

   PIN n_69725
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.482 0.0 106.51 0.163 ;
      END
   END n_69725

   PIN n_69742
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.346 0.0 23.374 0.163 ;
      END
   END n_69742

   PIN n_69765
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.034 0.0 106.062 0.163 ;
      END
   END n_69765

   PIN n_69846
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.226 0.0 98.254 0.163 ;
      END
   END n_69846

   PIN n_69856
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.218 0.0 23.246 0.163 ;
      END
   END n_69856

   PIN n_69945
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.89 0.0 11.918 0.163 ;
      END
   END n_69945

   PIN n_70024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.402 0.0 20.43 0.163 ;
      END
   END n_70024

   PIN n_70049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.634 0.0 11.662 0.163 ;
      END
   END n_70049

   PIN n_70182
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.874 0.0 101.902 0.163 ;
      END
   END n_70182

   PIN n_70208
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.954 0.0 11.982 0.163 ;
      END
   END n_70208

   PIN n_70223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.418 0.0 98.446 0.163 ;
      END
   END n_70223

   PIN n_70238
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.938 0.0 13.966 0.163 ;
      END
   END n_70238

   PIN n_70269
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.578 0.0 102.606 0.163 ;
      END
   END n_70269

   PIN n_70323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.578 0.0 102.606 0.163 ;
      END
   END n_70323

   PIN n_70327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.002 0.0 102.03 0.163 ;
      END
   END n_70327

   PIN n_70356
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.386 0.0 94.414 0.163 ;
      END
   END n_70356

   PIN n_70391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.29 0.0 98.318 0.163 ;
      END
   END n_70391

   PIN n_70403
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.354 0.0 106.382 0.082 ;
      END
   END n_70403

   PIN n_70473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.066 0.0 102.094 0.163 ;
      END
   END n_70473

   PIN n_70483
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.642 0.0 102.67 0.163 ;
      END
   END n_70483

   PIN n_70489
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.066 0.0 102.094 0.163 ;
      END
   END n_70489

   PIN n_70532
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.13 0.0 102.158 0.163 ;
      END
   END n_70532

   PIN n_70542
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.642 0.0 102.67 0.163 ;
      END
   END n_70542

   PIN n_70558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.914 0.0 20.942 0.163 ;
      END
   END n_70558

   PIN n_70643
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.146 0.0 100.174 0.163 ;
      END
   END n_70643

   PIN n_70646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.002 0.0 14.03 0.163 ;
      END
   END n_70646

   PIN n_70748
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.482 0.0 98.51 0.163 ;
      END
   END n_70748

   PIN n_70793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.162 0.0 98.19 0.163 ;
      END
   END n_70793

   PIN n_70794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.546 0.0 98.574 0.163 ;
      END
   END n_70794

   PIN n_70803
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.554 0.0 21.582 0.163 ;
      END
   END n_70803

   PIN n_70857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.834 0.0 94.862 0.163 ;
      END
   END n_70857

   PIN n_70928
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.61 0.0 98.638 0.163 ;
      END
   END n_70928

   PIN n_70933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.706 0.0 102.734 0.163 ;
      END
   END n_70933

   PIN n_71006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.77 0.0 102.798 0.163 ;
      END
   END n_71006

   PIN n_71030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.674 0.0 98.702 0.163 ;
      END
   END n_71030

   PIN n_71082
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.418 0.0 98.446 0.163 ;
      END
   END n_71082

   PIN n_71149
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.002 0.163 22.03 ;
      END
   END n_71149

   PIN n_71253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.802 0.163 18.83 ;
      END
   END n_71253

   PIN n_71285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.162 0.0 18.19 0.163 ;
      END
   END n_71285

   PIN n_71297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.074 0.0 25.102 0.163 ;
      END
   END n_71297

   PIN n_738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.874 0.0 5.902 0.163 ;
      END
   END n_738

   PIN n_75924
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.562 0.163 16.59 ;
      END
   END n_75924

   PIN n_75925
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.138 0.0 9.166 0.163 ;
      END
   END n_75925

   PIN n_76109
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.97 0.0 17.998 0.163 ;
      END
   END n_76109

   PIN n_76206
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.57 0.163 11.598 ;
      END
   END n_76206

   PIN n_76260
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.37 0.0 24.398 0.082 ;
      END
   END n_76260

   PIN n_76261
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.37 0.0 8.398 0.163 ;
      END
   END n_76261

   PIN n_76271
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.41 0.163 7.438 ;
      END
   END n_76271

   PIN n_76280
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.034 0.0 18.062 0.163 ;
      END
   END n_76280

   PIN n_76281
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.922 0.163 15.95 ;
      END
   END n_76281

   PIN n_76282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.786 0.163 12.814 ;
      END
   END n_76282

   PIN n_76283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.69 0.0 8.718 0.163 ;
      END
   END n_76283

   PIN n_76292
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.85 0.0 12.878 0.163 ;
      END
   END n_76292

   PIN n_76347
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.394 0.0 9.422 0.163 ;
      END
   END n_76347

   PIN n_76417
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.802 0.0 10.83 0.163 ;
      END
   END n_76417

   PIN n_76638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.626 0.0 8.654 0.163 ;
      END
   END n_76638

   PIN n_76852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.986 0.0 8.014 0.163 ;
      END
   END n_76852

   PIN n_76965
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.626 0.163 16.654 ;
      END
   END n_76965

   PIN n_77013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.778 0.0 9.806 0.163 ;
      END
   END n_77013

   PIN n_77047
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.114 0.0 8.142 0.163 ;
      END
   END n_77047

   PIN n_77053
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.274 0.163 20.302 ;
      END
   END n_77053

   PIN n_77442
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.986 0.0 8.014 0.163 ;
      END
   END n_77442

   PIN n_77600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.626 0.163 24.654 ;
      END
   END n_77600

   PIN n_78116
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.098 0.0 10.126 0.163 ;
      END
   END n_78116

   PIN n_823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.362 0.163 13.39 ;
      END
   END n_823

   PIN n_923
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.05 0.0 8.078 0.163 ;
      END
   END n_923

   PIN u0_L7_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.01 0.0 41.038 0.163 ;
      END
   END u0_L7_13_

   PIN u0_L7_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.85 0.0 44.878 0.163 ;
      END
   END u0_L7_3_

   PIN u0_L7_reg_14__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.746 0.0 37.774 0.163 ;
      END
   END u0_L7_reg_14__Q

   PIN u0_L7_reg_17__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.17 0.0 37.198 0.163 ;
      END
   END u0_L7_reg_17__Q

   PIN u0_L7_reg_18__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.114 0.0 88.142 0.163 ;
      END
   END u0_L7_reg_18__Q

   PIN u0_L8_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.154 0.0 63.182 0.163 ;
      END
   END u0_L8_12_

   PIN u0_L8_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.258 0.0 38.286 0.163 ;
      END
   END u0_L8_28_

   PIN u0_L8_reg_7__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.442 0.0 75.47 0.163 ;
      END
   END u0_L8_reg_7__Q

   PIN u0_L9_26_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.618 0.0 61.646 0.163 ;
      END
   END u0_L9_26_

   PIN u0_R10_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 175.581 3.506 175.744 3.534 ;
      END
   END u0_R10_23_

   PIN u0_R3_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.954 0.163 11.982 ;
      END
   END u0_R3_11_

   PIN u0_R4_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 19.954 0.163 19.982 ;
      END
   END u0_R4_1_

   PIN u0_R5_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.434 0.0 0.462 0.163 ;
      END
   END u0_R5_11_

   PIN u0_R5_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.178 0.0 8.206 0.163 ;
      END
   END u0_R5_14_

   PIN u0_R5_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.338 0.0 12.366 0.163 ;
      END
   END u0_R5_15_

   PIN u0_R5_19_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.938 0.0 5.966 0.163 ;
      END
   END u0_R5_19_

   PIN u0_R5_29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.338 0.0 44.366 0.163 ;
      END
   END u0_R5_29_

   PIN u0_R6_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.33 0.0 41.358 0.163 ;
      END
   END u0_R6_13_

   PIN u0_R6_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.042 0.0 13.07 0.163 ;
      END
   END u0_R6_1_

   PIN u0_R6_20_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.586 0.0 33.614 0.163 ;
      END
   END u0_R6_20_

   PIN u0_R6_30_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.066 0.0 30.094 0.163 ;
      END
   END u0_R6_30_

   PIN u0_R6_31_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.754 0.0 16.782 0.163 ;
      END
   END u0_R6_31_

   PIN u0_R6_32_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.818 0.0 16.846 0.163 ;
      END
   END u0_R6_32_

   PIN u0_R7_17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.674 0.0 18.702 0.163 ;
      END
   END u0_R7_17_

   PIN u0_R7_19_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.042 0.0 61.07 0.163 ;
      END
   END u0_R7_19_

   PIN u0_R7_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.89 0.0 35.918 0.163 ;
      END
   END u0_R7_7_

   PIN u0_R8_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.21 0.0 44.238 0.163 ;
      END
   END u0_R8_12_

   PIN u0_R8_17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.738 0.0 98.766 0.163 ;
      END
   END u0_R8_17_

   PIN u0_R8_20_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.674 0.0 26.702 0.163 ;
      END
   END u0_R8_20_

   PIN u0_R8_26_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.514 0.0 94.542 0.163 ;
      END
   END u0_R8_26_

   PIN u0_R8_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.186 0.0 83.214 0.163 ;
      END
   END u0_R8_3_

   PIN u0_R8_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.506 0.0 99.534 0.163 ;
      END
   END u0_R8_9_

   PIN u0_R9_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.786 0.0 140.814 0.163 ;
      END
   END u0_R9_12_

   PIN u0_R9_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.522 0.0 65.55 0.163 ;
      END
   END u0_R9_1_

   PIN u0_key_r_55_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.682 0.0 13.71 0.163 ;
      END
   END u0_key_r_55_

   PIN u0_uk_K_r_239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.01 0.0 25.038 0.163 ;
      END
   END u0_uk_K_r_239

   PIN u0_uk_K_r_264
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.45 0.163 6.478 ;
      END
   END u0_uk_K_r_264

   PIN u0_uk_K_r_349
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.746 0.0 13.774 0.163 ;
      END
   END u0_uk_K_r_349

   PIN u0_uk_K_r_353
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.93 0.0 2.958 0.163 ;
      END
   END u0_uk_K_r_353

   PIN u0_uk_K_r_361
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.298 0.0 5.326 0.163 ;
      END
   END u0_uk_K_r_361

   PIN u0_uk_K_r_373
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.642 0.163 6.67 ;
      END
   END u0_uk_K_r_373

   PIN u0_uk_K_r_383
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.666 0.0 7.694 0.163 ;
      END
   END u0_uk_K_r_383

   PIN u0_uk_K_r_387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.058 0.163 11.086 ;
      END
   END u0_uk_K_r_387

   PIN u0_uk_K_r_390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.818 0.163 8.846 ;
      END
   END u0_uk_K_r_390

   PIN u0_uk_K_r_399
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.498 0.163 8.526 ;
      END
   END u0_uk_K_r_399

   PIN u0_uk_K_r_412
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.698 0.0 11.726 0.163 ;
      END
   END u0_uk_K_r_412

   PIN u0_uk_K_r_433
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.082 0.0 4.11 0.163 ;
      END
   END u0_uk_K_r_433

   PIN u0_uk_K_r_436
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.106 0.0 5.134 0.163 ;
      END
   END u0_uk_K_r_436

   PIN u0_uk_K_r_463
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.018 0.163 12.046 ;
      END
   END u0_uk_K_r_463

   PIN u0_uk_K_r_469
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.442 0.0 3.47 0.163 ;
      END
   END u0_uk_K_r_469

   PIN u0_uk_K_r_492
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.826 0.0 3.854 0.163 ;
      END
   END u0_uk_K_r_492

   PIN u0_uk_K_r_518
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.114 0.0 8.142 0.163 ;
      END
   END u0_uk_K_r_518

   PIN u0_uk_K_r_523
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.69 0.163 16.718 ;
      END
   END u0_uk_K_r_523

   PIN u0_uk_K_r_547
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.658 0.0 4.686 0.163 ;
      END
   END u0_uk_K_r_547

   PIN u1_IP_22_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.434 0.0 24.462 0.163 ;
      END
   END u1_IP_22_

   PIN u1_L11_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.13 0.0 102.158 0.163 ;
      END
   END u1_L11_7_

   PIN u1_R10_29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.042 0.163 13.07 ;
      END
   END u1_R10_29_

   PIN u1_R10_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.794 0.163 7.822 ;
      END
   END u1_R10_4_

   PIN u1_desIn_r_reg_28__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.426 0.0 29.454 0.163 ;
      END
   END u1_desIn_r_reg_28__Q

   PIN u1_desIn_r_reg_54__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.546 0.0 18.574 0.163 ;
      END
   END u1_desIn_r_reg_54__Q

   PIN u2_L7_reg_12__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.426 0.0 125.454 0.163 ;
      END
   END u2_L7_reg_12__Q

   PIN u2_L7_reg_7__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.362 0.0 117.39 0.163 ;
      END
   END u2_L7_reg_7__Q

   PIN FE_OFN1018_n_6197
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.018 0.0 12.046 0.163 ;
      END
   END FE_OFN1018_n_6197

   PIN FE_OFN1021_n_3701
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.074 0.0 1.102 0.163 ;
      END
   END FE_OFN1021_n_3701

   PIN FE_OFN1068_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.946 0.0 8.974 0.163 ;
      END
   END FE_OFN1068_n_116

   PIN FE_OFN1094_g303299_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.458 0.0 1.486 0.163 ;
      END
   END FE_OFN1094_g303299_p

   PIN FE_OFN1105_n_6021
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.93 0.0 18.958 0.163 ;
      END
   END FE_OFN1105_n_6021

   PIN FE_OFN1224_n_6583
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.802 0.0 26.83 0.163 ;
      END
   END FE_OFN1224_n_6583

   PIN FE_OFN1292_n_4098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.602 0.0 7.63 0.163 ;
      END
   END FE_OFN1292_n_4098

   PIN FE_OFN1338_n_117596
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.794 0.0 63.822 0.163 ;
      END
   END FE_OFN1338_n_117596

   PIN FE_OFN1381_n_6875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.058 0.0 51.086 0.163 ;
      END
   END FE_OFN1381_n_6875

   PIN FE_OFN1578_n_3047
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.162 0.0 2.19 0.163 ;
      END
   END FE_OFN1578_n_3047

   PIN FE_OFN1646_n_6731
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.066 0.0 54.094 0.163 ;
      END
   END FE_OFN1646_n_6731

   PIN FE_OFN1735_n_64033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 28.338 0.082 28.366 ;
      END
   END FE_OFN1735_n_64033

   PIN FE_OFN1933_n_69492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.882 0.0 24.91 0.163 ;
      END
   END FE_OFN1933_n_69492

   PIN FE_OFN1958_n_6873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.258 0.0 30.286 0.163 ;
      END
   END FE_OFN1958_n_6873

   PIN FE_OFN2009_n_27918
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.418 0.0 18.446 0.163 ;
      END
   END FE_OFN2009_n_27918

   PIN FE_OFN2013_n_23906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.954 0.0 3.982 0.163 ;
      END
   END FE_OFN2013_n_23906

   PIN FE_OFN2114_n_19614
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.098 0.0 18.126 0.163 ;
      END
   END FE_OFN2114_n_19614

   PIN FE_OFN2221_g302057_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.946 0.0 0.974 0.163 ;
      END
   END FE_OFN2221_g302057_p

   PIN FE_OFN2276_n_27867
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.122 0.0 11.15 0.163 ;
      END
   END FE_OFN2276_n_27867

   PIN FE_OFN2316_n_65154
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.722 0.0 20.75 0.163 ;
      END
   END FE_OFN2316_n_65154

   PIN FE_OFN2333_n_23919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.57 0.163 3.598 ;
      END
   END FE_OFN2333_n_23919

   PIN FE_OFN2351_n_27890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.754 0.0 8.782 0.163 ;
      END
   END FE_OFN2351_n_27890

   PIN FE_OFN2406_n_13312
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.498 0.0 0.526 0.163 ;
      END
   END FE_OFN2406_n_13312

   PIN FE_OFN2417_n_26365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.026 0.163 55.054 ;
      END
   END FE_OFN2417_n_26365

   PIN FE_OFN2472_n_117820
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.874 0.0 5.902 0.163 ;
      END
   END FE_OFN2472_n_117820

   PIN FE_OFN2503_n_5437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.69 0.0 24.718 0.163 ;
      END
   END FE_OFN2503_n_5437

   PIN FE_OFN2504_n_4918
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.546 0.0 2.574 0.163 ;
      END
   END FE_OFN2504_n_4918

   PIN FE_OFN2537_n_65517
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.482 0.0 2.51 0.163 ;
      END
   END FE_OFN2537_n_65517

   PIN FE_OFN2677_n_23958
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.554 0.0 13.582 0.163 ;
      END
   END FE_OFN2677_n_23958

   PIN FE_OFN2719_n_25980
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.05 0.0 8.078 0.163 ;
      END
   END FE_OFN2719_n_25980

   PIN FE_OFN2786_n_5684
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.762 0.0 11.79 0.163 ;
      END
   END FE_OFN2786_n_5684

   PIN FE_OFN2930_n_4064
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.042 0.0 5.07 0.163 ;
      END
   END FE_OFN2930_n_4064

   PIN FE_OFN2965_n_4653
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.066 0.0 6.094 0.163 ;
      END
   END FE_OFN2965_n_4653

   PIN FE_OFN2975_n_65768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.01 0.0 1.038 0.163 ;
      END
   END FE_OFN2975_n_65768

   PIN FE_OFN2982_n_65436
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.002 0.0 14.03 0.163 ;
      END
   END FE_OFN2982_n_65436

   PIN FE_OFN2993_n_6198
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.85 0.0 4.878 0.163 ;
      END
   END FE_OFN2993_n_6198

   PIN FE_OFN3017_n_69766
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.202 0.0 25.23 0.163 ;
      END
   END FE_OFN3017_n_69766

   PIN FE_OFN3049_n_3016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.69 0.0 8.718 0.163 ;
      END
   END FE_OFN3049_n_3016

   PIN FE_OFN3146_n_35477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.482 0.0 90.51 0.163 ;
      END
   END FE_OFN3146_n_35477

   PIN FE_OFN3152_n_25832
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.634 0.0 11.662 0.163 ;
      END
   END FE_OFN3152_n_25832

   PIN FE_OFN3164_n_2780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.666 0.0 7.694 0.163 ;
      END
   END FE_OFN3164_n_2780

   PIN FE_OFN3226_g302039_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.466 0.0 4.494 0.163 ;
      END
   END FE_OFN3226_g302039_p

   PIN FE_OFN3240_n_4790
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.434 0.163 8.462 ;
      END
   END FE_OFN3240_n_4790

   PIN FE_OFN324_n_70684
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.354 0.0 106.382 0.163 ;
      END
   END FE_OFN324_n_70684

   PIN FE_OFN326_n_70685
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.386 0.0 102.414 0.163 ;
      END
   END FE_OFN326_n_70685

   PIN FE_OFN3278_n_39
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.202 0.0 1.23 0.163 ;
      END
   END FE_OFN3278_n_39

   PIN FE_OFN3318_n_500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.666 94.638 31.694 94.72 ;
      END
   END FE_OFN3318_n_500

   PIN FE_OFN3319_n_500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.642 0.082 30.67 ;
      END
   END FE_OFN3319_n_500

   PIN FE_OFN3365_n_5443
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.386 0.0 6.414 0.163 ;
      END
   END FE_OFN3365_n_5443

   PIN FE_OFN3399_n_7096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.162 0.0 2.19 0.163 ;
      END
   END FE_OFN3399_n_7096

   PIN FE_OFN3463_n_67106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.298 0.163 13.326 ;
      END
   END FE_OFN3463_n_67106

   PIN FE_OFN3485_n_1596
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.634 0.0 3.662 0.163 ;
      END
   END FE_OFN3485_n_1596

   PIN FE_OFN3516_n_23820
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.258 0.163 6.286 ;
      END
   END FE_OFN3516_n_23820

   PIN FE_OFN3542_g302047_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.842 0.0 1.87 0.163 ;
      END
   END FE_OFN3542_g302047_p

   PIN FE_OFN3627_n_4557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.738 0.0 10.766 0.163 ;
      END
   END FE_OFN3627_n_4557

   PIN FE_OFN373_n_66358
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.89 0.0 11.918 0.163 ;
      END
   END FE_OFN373_n_66358

   PIN FE_OFN375_n_65823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.154 0.0 7.182 0.163 ;
      END
   END FE_OFN375_n_65823

   PIN FE_OFN3784_n_60
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.626 0.163 8.654 ;
      END
   END FE_OFN3784_n_60

   PIN FE_OFN3799_n_23840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.17 0.163 5.198 ;
      END
   END FE_OFN3799_n_23840

   PIN FE_OFN3858_n_68782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.01 0.0 17.038 0.163 ;
      END
   END FE_OFN3858_n_68782

   PIN FE_OFN3909_n_5532
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.722 0.0 4.75 0.163 ;
      END
   END FE_OFN3909_n_5532

   PIN FE_OFN3914_n_29934
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.954 0.0 115.982 0.163 ;
      END
   END FE_OFN3914_n_29934

   PIN FE_OFN3965_n_9884
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.866 0.163 10.894 ;
      END
   END FE_OFN3965_n_9884

   PIN FE_OFN4124_g302043_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.522 0.0 1.55 0.163 ;
      END
   END FE_OFN4124_g302043_p

   PIN FE_OFN4143_n_29936
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.914 0.0 44.942 0.163 ;
      END
   END FE_OFN4143_n_29936

   PIN FE_OFN4244_n_29500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.946 0.0 56.974 0.163 ;
      END
   END FE_OFN4244_n_29500

   PIN FE_OFN4315_n_104
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.418 0.0 10.446 0.082 ;
      END
   END FE_OFN4315_n_104

   PIN FE_OFN4359_n_20
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.41 0.0 7.438 0.082 ;
      END
   END FE_OFN4359_n_20

   PIN FE_OFN4412_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.73 0.082 7.758 ;
      END
   END FE_OFN4412_decrypt

   PIN FE_OFN4422_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.714 0.082 9.742 ;
      END
   END FE_OFN4422_decrypt

   PIN FE_OFN4476_n_39
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.746 0.0 5.774 0.082 ;
      END
   END FE_OFN4476_n_39

   PIN FE_OFN4517_n_13659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.674 0.0 10.702 0.163 ;
      END
   END FE_OFN4517_n_13659

   PIN FE_OFN4612_n_201
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.202 0.0 1.23 0.163 ;
      END
   END FE_OFN4612_n_201

   PIN FE_OFN4797_n_21953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.514 0.163 6.542 ;
      END
   END FE_OFN4797_n_21953

   PIN FE_OFN663_n_32304
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.882 0.0 48.91 0.163 ;
      END
   END FE_OFN663_n_32304

   PIN FE_OFN669_n_32833
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.122 0.0 75.15 0.163 ;
      END
   END FE_OFN669_n_32833

   PIN FE_OFN677_n_30310
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.09 0.0 119.118 0.163 ;
      END
   END FE_OFN677_n_30310

   PIN FE_OFN683_n_117971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.186 0.163 51.214 ;
      END
   END FE_OFN683_n_117971

   PIN FE_OFN692_n_27625
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.962 0.163 54.99 ;
      END
   END FE_OFN692_n_27625

   PIN FE_OFN852_n_3353
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.89 0.0 3.918 0.163 ;
      END
   END FE_OFN852_n_3353

   PIN FE_OFN910_n_21872
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.322 0.163 6.35 ;
      END
   END FE_OFN910_n_21872

   PIN FE_OFN947_n_3795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.754 0.163 8.782 ;
      END
   END FE_OFN947_n_3795

   PIN FE_OFN972_n_63299
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.106 0.163 5.134 ;
      END
   END FE_OFN972_n_63299

   PIN g205805_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.354 0.0 74.382 0.163 ;
      END
   END g205805_sb

   PIN g231413_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.37 0.163 24.398 ;
      END
   END g231413_p

   PIN g233023_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.09 94.557 23.118 94.72 ;
      END
   END g233023_p

   PIN g233195_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.898 0.0 6.926 0.163 ;
      END
   END g233195_p

   PIN g235329_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.746 0.0 21.774 0.163 ;
      END
   END g235329_p

   PIN g265215_p2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.37 0.0 88.398 0.163 ;
      END
   END g265215_p2

   PIN g266100_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.346 0.0 63.374 0.163 ;
      END
   END g266100_p

   PIN g267780_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.538 0.0 71.566 0.163 ;
      END
   END g267780_p

   PIN g267919_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.506 0.0 75.534 0.163 ;
      END
   END g267919_p

   PIN g268186_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.106 0.0 69.134 0.163 ;
      END
   END g268186_p

   PIN g268308_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.458 0.0 65.486 0.163 ;
      END
   END g268308_p

   PIN g268393_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.818 0.0 48.846 0.163 ;
      END
   END g268393_p

   PIN g268990_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.818 0.0 40.846 0.163 ;
      END
   END g268990_p

   PIN g269848_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.674 0.0 114.702 0.163 ;
      END
   END g269848_p

   PIN g270852_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.386 0.0 62.414 0.163 ;
      END
   END g270852_p

   PIN g271549_p1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.194 0.0 62.222 0.163 ;
      END
   END g271549_p1

   PIN g271686_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.882 0.0 56.91 0.163 ;
      END
   END g271686_p

   PIN g271749_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.354 0.0 58.382 0.163 ;
      END
   END g271749_p

   PIN g271784_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.186 0.0 59.214 0.163 ;
      END
   END g271784_p

   PIN g271972_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.45 0.0 62.478 0.163 ;
      END
   END g271972_p

   PIN g272788_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.266 0.0 57.294 0.163 ;
      END
   END g272788_p

   PIN g272818_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.722 0.0 12.75 0.163 ;
      END
   END g272818_sb

   PIN g272848_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.274 0.0 12.302 0.163 ;
      END
   END g272848_p

   PIN g273938_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.242 0.163 8.27 ;
      END
   END g273938_p

   PIN g273953_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.554 0.163 13.582 ;
      END
   END g273953_p

   PIN g278067_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.338 0.0 4.366 0.163 ;
      END
   END g278067_p

   PIN g279539_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.514 0.0 6.542 0.163 ;
      END
   END g279539_db

   PIN g279539_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.57 0.0 3.598 0.163 ;
      END
   END g279539_sb

   PIN g302013_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.578 0.163 6.606 ;
      END
   END g302013_p

   PIN g302028_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.01 0.0 1.038 0.163 ;
      END
   END g302028_p

   PIN g302042_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.754 0.163 16.782 ;
      END
   END g302042_p

   PIN g302689_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.642 0.163 6.67 ;
      END
   END g302689_p

   PIN g303333_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.69 0.163 8.718 ;
      END
   END g303333_p

   PIN g303373_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.842 0.0 1.87 0.163 ;
      END
   END g303373_p

   PIN g304261_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.882 0.0 0.91 0.163 ;
      END
   END g304261_p

   PIN g304290_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.778 0.0 1.806 0.163 ;
      END
   END g304290_p

   PIN g304292_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.29 0.0 2.318 0.163 ;
      END
   END g304292_p

   PIN g305157_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.13 0.0 30.158 0.163 ;
      END
   END g305157_p

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.234 0.0 13.262 0.163 ;
      END
   END ispd_clk

   PIN key1_19_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.546 94.557 2.574 94.72 ;
      END
   END key1_19_

   PIN key1_55_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.426 94.557 29.454 94.72 ;
      END
   END key1_55_

   PIN key3_19_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.826 94.557 3.854 94.72 ;
      END
   END key3_19_

   PIN key3_55_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.266 94.557 33.294 94.72 ;
      END
   END key3_55_

   PIN n_1023
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END n_1023

   PIN n_10608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.914 0.0 4.942 0.163 ;
      END
   END n_10608

   PIN n_108553
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.626 0.0 40.654 0.163 ;
      END
   END n_108553

   PIN n_108562
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.346 0.163 15.374 ;
      END
   END n_108562

   PIN n_108697
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.658 0.163 20.686 ;
      END
   END n_108697

   PIN n_108698
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.426 0.0 29.454 0.163 ;
      END
   END n_108698

   PIN n_108729
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.914 0.163 12.942 ;
      END
   END n_108729

   PIN n_108760
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.17 0.0 13.198 0.163 ;
      END
   END n_108760

   PIN n_108971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.594 0.0 4.622 0.163 ;
      END
   END n_108971

   PIN n_109090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.13 0.0 110.158 0.163 ;
      END
   END n_109090

   PIN n_109137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.978 0.0 13.006 0.163 ;
      END
   END n_109137

   PIN n_109138
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.106 0.0 13.134 0.163 ;
      END
   END n_109138

   PIN n_112756
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.074 94.557 41.102 94.72 ;
      END
   END n_112756

   PIN n_112757
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.01 94.557 41.038 94.72 ;
      END
   END n_112757

   PIN n_112829
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.722 0.0 44.75 0.163 ;
      END
   END n_112829

   PIN n_116914
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.714 0.0 9.742 0.163 ;
      END
   END n_116914

   PIN n_116948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.562 0.0 16.59 0.163 ;
      END
   END n_116948

   PIN n_117298
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.106 0.0 53.134 0.163 ;
      END
   END n_117298

   PIN n_117339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.81 0.0 5.838 0.163 ;
      END
   END n_117339

   PIN n_117340
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.818 0.163 16.846 ;
      END
   END n_117340

   PIN n_117465
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.786 0.0 12.814 0.163 ;
      END
   END n_117465

   PIN n_117466
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.834 0.0 6.862 0.163 ;
      END
   END n_117466

   PIN n_117596
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.73 0.0 71.758 0.163 ;
      END
   END n_117596

   PIN n_117600
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.418 0.0 66.446 0.163 ;
      END
   END n_117600

   PIN n_117902
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.01 0.163 9.038 ;
      END
   END n_117902

   PIN n_118304
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.81 0.0 45.838 0.163 ;
      END
   END n_118304

   PIN n_118305
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.618 0.0 45.646 0.163 ;
      END
   END n_118305

   PIN n_118591
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.298 94.557 5.326 94.72 ;
      END
   END n_118591

   PIN n_118596
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.674 0.0 2.702 0.163 ;
      END
   END n_118596

   PIN n_118598
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.746 94.557 5.774 94.72 ;
      END
   END n_118598

   PIN n_1263
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.234 0.0 5.262 0.163 ;
      END
   END n_1263

   PIN n_1266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.274 0.0 4.302 0.163 ;
      END
   END n_1266

   PIN n_1281
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.042 0.163 5.07 ;
      END
   END n_1281

   PIN n_1387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.074 0.0 9.102 0.163 ;
      END
   END n_1387

   PIN n_13938
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.978 0.0 5.006 0.163 ;
      END
   END n_13938

   PIN n_1489
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END n_1489

   PIN n_1501
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.914 0.0 4.942 0.163 ;
      END
   END n_1501

   PIN n_1504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.89 0.0 3.918 0.163 ;
      END
   END n_1504

   PIN n_1529
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.714 0.0 1.742 0.163 ;
      END
   END n_1529

   PIN n_155186
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.882 0.0 40.91 0.163 ;
      END
   END n_155186

   PIN n_1593
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.802 0.163 10.83 ;
      END
   END n_1593

   PIN n_1646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.506 0.163 3.534 ;
      END
   END n_1646

   PIN n_18158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.09 0.163 7.118 ;
      END
   END n_18158

   PIN n_18380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.946 0.0 0.974 0.163 ;
      END
   END n_18380

   PIN n_18386
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.97 0.163 9.998 ;
      END
   END n_18386

   PIN n_1848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.858 0.0 7.886 0.163 ;
      END
   END n_1848

   PIN n_18639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.826 0.0 3.854 0.163 ;
      END
   END n_18639

   PIN n_18670
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.898 0.0 6.926 0.163 ;
      END
   END n_18670

   PIN n_18679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.322 0.163 70.35 ;
      END
   END n_18679

   PIN n_1878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.97 0.0 1.998 0.163 ;
      END
   END n_1878

   PIN n_18862
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.706 0.163 6.734 ;
      END
   END n_18862

   PIN n_19056
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.882 0.0 0.91 0.163 ;
      END
   END n_19056

   PIN n_19424
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.458 0.0 1.486 0.163 ;
      END
   END n_19424

   PIN n_19436
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.186 0.163 11.214 ;
      END
   END n_19436

   PIN n_19692
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.69 0.163 8.718 ;
      END
   END n_19692

   PIN n_19693
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.978 0.163 5.006 ;
      END
   END n_19693

   PIN n_19844
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.546 0.163 66.574 ;
      END
   END n_19844

   PIN n_19868
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.906 0.0 1.934 0.163 ;
      END
   END n_19868

   PIN n_20239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.266 0.163 9.294 ;
      END
   END n_20239

   PIN n_20284
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.482 0.163 66.51 ;
      END
   END n_20284

   PIN n_20529
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.914 0.163 4.942 ;
      END
   END n_20529

   PIN n_20542
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.85 0.163 4.878 ;
      END
   END n_20542

   PIN n_20744
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.394 0.0 1.422 0.163 ;
      END
   END n_20744

   PIN n_20818
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.386 0.163 6.414 ;
      END
   END n_20818

   PIN n_21311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.594 0.0 4.622 0.163 ;
      END
   END n_21311

   PIN n_2155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.586 0.0 1.614 0.163 ;
      END
   END n_2155

   PIN n_21823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.506 0.163 11.534 ;
      END
   END n_21823

   PIN n_21905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.77 0.163 6.798 ;
      END
   END n_21905

   PIN n_21912
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.434 0.0 8.462 0.163 ;
      END
   END n_21912

   PIN n_21921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.874 0.163 77.902 ;
      END
   END n_21921

   PIN n_21949
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.89 0.163 19.918 ;
      END
   END n_21949

   PIN n_21999
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.026 0.0 7.054 0.163 ;
      END
   END n_21999

   PIN n_22036
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.306 0.163 16.334 ;
      END
   END n_22036

   PIN n_22173
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.73 0.0 7.758 0.163 ;
      END
   END n_22173

   PIN n_22174
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.45 0.0 6.478 0.163 ;
      END
   END n_22174

   PIN n_22255
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.45 0.0 6.478 0.163 ;
      END
   END n_22255

   PIN n_22325
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.794 0.0 7.822 0.163 ;
      END
   END n_22325

   PIN n_22338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.17 0.0 13.198 0.163 ;
      END
   END n_22338

   PIN n_22350
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.682 0.0 5.71 0.163 ;
      END
   END n_22350

   PIN n_22352
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.106 0.0 5.134 0.163 ;
      END
   END n_22352

   PIN n_22359
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.09 0.0 7.118 0.163 ;
      END
   END n_22359

   PIN n_22392
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.562 0.0 0.59 0.163 ;
      END
   END n_22392

   PIN n_22454
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.882 0.163 16.91 ;
      END
   END n_22454

   PIN n_22603
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.586 0.163 9.614 ;
      END
   END n_22603

   PIN n_22612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.842 0.163 9.87 ;
      END
   END n_22612

   PIN n_22800
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.786 0.0 4.814 0.163 ;
      END
   END n_22800

   PIN n_22836
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.85 0.163 12.878 ;
      END
   END n_22836

   PIN n_22929
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.914 0.163 12.942 ;
      END
   END n_22929

   PIN n_22932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.13 0.0 6.158 0.163 ;
      END
   END n_22932

   PIN n_22937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.634 0.163 11.662 ;
      END
   END n_22937

   PIN n_23053
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.538 0.0 7.566 0.163 ;
      END
   END n_23053

   PIN n_23062
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.53 0.0 4.558 0.163 ;
      END
   END n_23062

   PIN n_23073
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.258 0.0 6.286 0.163 ;
      END
   END n_23073

   PIN n_23091
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.642 0.0 6.67 0.163 ;
      END
   END n_23091

   PIN n_23165
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.946 0.163 16.974 ;
      END
   END n_23165

   PIN n_23219
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.498 0.163 8.526 ;
      END
   END n_23219

   PIN n_2332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.706 0.0 6.734 0.163 ;
      END
   END n_2332

   PIN n_2334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.722 0.163 20.75 ;
      END
   END n_2334

   PIN n_23606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.218 0.0 7.246 0.163 ;
      END
   END n_23606

   PIN n_23635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.258 0.0 6.286 0.163 ;
      END
   END n_23635

   PIN n_23694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.626 0.0 8.654 0.163 ;
      END
   END n_23694

   PIN n_23721
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.562 0.0 8.59 0.163 ;
      END
   END n_23721

   PIN n_23876
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.834 0.163 6.862 ;
      END
   END n_23876

   PIN n_24030
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.898 0.163 6.926 ;
      END
   END n_24030

   PIN n_24048
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.378 0.163 3.406 ;
      END
   END n_24048

   PIN n_2435
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.786 0.163 4.814 ;
      END
   END n_2435

   PIN n_24781
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.722 0.163 4.75 ;
      END
   END n_24781

   PIN n_2483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.234 0.0 5.262 0.163 ;
      END
   END n_2483

   PIN n_2504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.034 0.0 2.062 0.163 ;
      END
   END n_2504

   PIN n_25070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.146 0.163 4.174 ;
      END
   END n_25070

   PIN n_25088
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.97 94.557 17.998 94.72 ;
      END
   END n_25088

   PIN n_25090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.066 94.557 14.094 94.72 ;
      END
   END n_25090

   PIN n_25102
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.138 94.557 1.166 94.72 ;
      END
   END n_25102

   PIN n_25130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.818 94.557 0.846 94.72 ;
      END
   END n_25130

   PIN n_25224
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.474 0.163 7.502 ;
      END
   END n_25224

   PIN n_25227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.658 0.163 4.686 ;
      END
   END n_25227

   PIN n_25228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.946 0.163 8.974 ;
      END
   END n_25228

   PIN n_25317
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.41 0.163 7.438 ;
      END
   END n_25317

   PIN n_25375
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.594 0.163 4.622 ;
      END
   END n_25375

   PIN n_25412
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.346 0.163 7.374 ;
      END
   END n_25412

   PIN n_2549
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.658 0.0 12.686 0.163 ;
      END
   END n_2549

   PIN n_25591
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.13 94.557 14.158 94.72 ;
      END
   END n_25591

   PIN n_25662
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.082 0.163 20.11 ;
      END
   END n_25662

   PIN n_25669
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.066 94.557 14.094 94.72 ;
      END
   END n_25669

   PIN n_25671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.842 94.557 17.87 94.72 ;
      END
   END n_25671

   PIN n_25677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.002 94.557 14.03 94.72 ;
      END
   END n_25677

   PIN n_25679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.362 94.557 5.39 94.72 ;
      END
   END n_25679

   PIN n_25713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.842 94.557 17.87 94.72 ;
      END
   END n_25713

   PIN n_25727
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.178 0.163 24.206 ;
      END
   END n_25727

   PIN n_25764
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.306 0.163 24.334 ;
      END
   END n_25764

   PIN n_25771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.018 0.163 4.046 ;
      END
   END n_25771

   PIN n_25794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.97 0.0 1.998 0.163 ;
      END
   END n_25794

   PIN n_25810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.722 0.0 36.75 0.163 ;
      END
   END n_25810

   PIN n_25823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.13 0.163 14.158 ;
      END
   END n_25823

   PIN n_25837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.978 0.0 29.006 0.163 ;
      END
   END n_25837

   PIN n_25849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.146 0.0 12.174 0.163 ;
      END
   END n_25849

   PIN n_25856
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.322 0.0 6.35 0.163 ;
      END
   END n_25856

   PIN n_25870
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.242 0.0 8.27 0.163 ;
      END
   END n_25870

   PIN n_25888
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.29 0.0 10.318 0.163 ;
      END
   END n_25888

   PIN n_25889
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.986 0.163 8.014 ;
      END
   END n_25889

   PIN n_25895
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.434 0.163 8.462 ;
      END
   END n_25895

   PIN n_25935
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.57 0.0 59.598 0.163 ;
      END
   END n_25935

   PIN n_26069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.962 0.0 14.99 0.163 ;
      END
   END n_26069

   PIN n_26071
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.194 0.163 14.222 ;
      END
   END n_26071

   PIN n_26153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 94.557 25.614 94.72 ;
      END
   END n_26153

   PIN n_26374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.858 0.163 7.886 ;
      END
   END n_26374

   PIN n_26377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.058 0.163 3.086 ;
      END
   END n_26377

   PIN n_26491
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.17 0.0 29.198 0.163 ;
      END
   END n_26491

   PIN n_26510
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.714 0.0 17.742 0.163 ;
      END
   END n_26510

   PIN n_26547
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.682 0.082 13.71 ;
      END
   END n_26547

   PIN n_26553
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.05 0.163 16.078 ;
      END
   END n_26553

   PIN n_26558
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.226 0.0 2.254 0.163 ;
      END
   END n_26558

   PIN n_26622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.282 0.163 15.31 ;
      END
   END n_26622

   PIN n_2663
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.138 0.0 25.166 0.163 ;
      END
   END n_2663

   PIN n_26632
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 13.298 0.163 13.326 ;
      END
   END n_26632

   PIN n_26638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.802 0.163 2.83 ;
      END
   END n_26638

   PIN n_26672
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.386 0.163 14.414 ;
      END
   END n_26672

   PIN n_26763
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.002 0.163 14.03 ;
      END
   END n_26763

   PIN n_26765
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.322 0.163 14.35 ;
      END
   END n_26765

   PIN n_26785
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.874 0.163 13.902 ;
      END
   END n_26785

   PIN n_2679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.274 0.163 4.302 ;
      END
   END n_2679

   PIN n_26983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.978 0.163 13.006 ;
      END
   END n_26983

   PIN n_27075
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.426 0.163 13.454 ;
      END
   END n_27075

   PIN n_2708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.562 0.163 8.59 ;
      END
   END n_2708

   PIN n_27099
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.266 0.0 1.294 0.163 ;
      END
   END n_27099

   PIN n_27127
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.866 0.163 2.894 ;
      END
   END n_27127

   PIN n_27563
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.834 0.163 6.862 ;
      END
   END n_27563

   PIN n_27603
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.954 0.163 27.982 ;
      END
   END n_27603

   PIN n_27616
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.922 0.0 7.95 0.163 ;
      END
   END n_27616

   PIN n_27646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.338 0.163 20.366 ;
      END
   END n_27646

   PIN n_27654
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.914 0.0 28.942 0.163 ;
      END
   END n_27654

   PIN n_27671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.226 0.163 74.254 ;
      END
   END n_27671

   PIN n_27702
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.386 0.163 70.414 ;
      END
   END n_27702

   PIN n_27743
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.338 0.163 12.366 ;
      END
   END n_27743

   PIN n_27794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.57 0.0 11.598 0.163 ;
      END
   END n_27794

   PIN n_2780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.53 0.163 4.558 ;
      END
   END n_2780

   PIN n_27806
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.506 0.0 11.534 0.163 ;
      END
   END n_27806

   PIN n_27815
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.802 0.0 18.83 0.163 ;
      END
   END n_27815

   PIN n_27847
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.002 0.0 6.03 0.163 ;
      END
   END n_27847

   PIN n_27858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.194 0.0 102.222 0.163 ;
      END
   END n_27858

   PIN n_27869
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.186 0.0 83.214 0.163 ;
      END
   END n_27869

   PIN n_27978
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.01 0.0 33.038 0.163 ;
      END
   END n_27978

   PIN n_27984
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.138 0.0 33.166 0.163 ;
      END
   END n_27984

   PIN n_28031
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.37 0.0 32.398 0.163 ;
      END
   END n_28031

   PIN n_28036
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.65 0.0 33.678 0.163 ;
      END
   END n_28036

   PIN n_28044
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.794 0.0 31.822 0.163 ;
      END
   END n_28044

   PIN n_28072
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.69 0.0 32.718 0.163 ;
      END
   END n_28072

   PIN n_281
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.442 0.163 3.47 ;
      END
   END n_281

   PIN n_28101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.786 0.0 36.814 0.163 ;
      END
   END n_28101

   PIN n_28135
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.53 0.0 52.558 0.163 ;
      END
   END n_28135

   PIN n_28136
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.338 0.0 52.366 0.163 ;
      END
   END n_28136

   PIN n_28138
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.882 0.0 56.91 0.163 ;
      END
   END n_28138

   PIN n_28140
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.714 0.0 57.742 0.163 ;
      END
   END n_28140

   PIN n_28166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.722 0.0 12.75 0.163 ;
      END
   END n_28166

   PIN n_28204
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.986 0.0 56.014 0.163 ;
      END
   END n_28204

   PIN n_28212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.618 0.0 29.646 0.163 ;
      END
   END n_28212

   PIN n_28230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.29 0.0 34.318 0.163 ;
      END
   END n_28230

   PIN n_28237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.882 0.0 32.91 0.082 ;
      END
   END n_28237

   PIN n_28309
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.754 0.0 32.782 0.082 ;
      END
   END n_28309

   PIN n_28396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.978 0.0 61.006 0.163 ;
      END
   END n_28396

   PIN n_28398
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.714 0.0 33.742 0.163 ;
      END
   END n_28398

   PIN n_28447
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.202 0.0 33.23 0.163 ;
      END
   END n_28447

   PIN n_28448
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.738 0.0 58.766 0.163 ;
      END
   END n_28448

   PIN n_28501
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.106 0.0 37.134 0.163 ;
      END
   END n_28501

   PIN n_28504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.562 0.0 32.59 0.163 ;
      END
   END n_28504

   PIN n_28534
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.914 0.0 36.942 0.163 ;
      END
   END n_28534

   PIN n_28606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.626 0.0 32.654 0.163 ;
      END
   END n_28606

   PIN n_28621
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.722 0.0 36.75 0.163 ;
      END
   END n_28621

   PIN n_28622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.77 0.0 30.798 0.163 ;
      END
   END n_28622

   PIN n_28639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.674 0.0 58.702 0.163 ;
      END
   END n_28639

   PIN n_28712
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.33 0.0 33.358 0.163 ;
      END
   END n_28712

   PIN n_28713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.114 0.0 32.142 0.163 ;
      END
   END n_28713

   PIN n_28715
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.73 0.0 31.758 0.163 ;
      END
   END n_28715

   PIN n_28717
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.346 0.0 31.374 0.163 ;
      END
   END n_28717

   PIN n_28780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.042 0.0 37.07 0.163 ;
      END
   END n_28780

   PIN n_28805
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.658 0.0 36.686 0.163 ;
      END
   END n_28805

   PIN n_28859
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.882 0.0 32.91 0.163 ;
      END
   END n_28859

   PIN n_2887
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.018 0.163 20.046 ;
      END
   END n_2887

   PIN n_28880
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.746 0.0 61.774 0.163 ;
      END
   END n_28880

   PIN n_29030
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.954 0.0 59.982 0.163 ;
      END
   END n_29030

   PIN n_29061
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.002 0.0 30.03 0.163 ;
      END
   END n_29061

   PIN n_29110
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.562 0.0 56.59 0.163 ;
      END
   END n_29110

   PIN n_29123
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.602 0.0 31.63 0.163 ;
      END
   END n_29123

   PIN n_29127
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.53 0.0 36.558 0.163 ;
      END
   END n_29127

   PIN n_29141
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.29 0.0 58.318 0.163 ;
      END
   END n_29141

   PIN n_29150
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.386 0.0 62.414 0.163 ;
      END
   END n_29150

   PIN n_29151
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.442 0.0 59.47 0.163 ;
      END
   END n_29151

   PIN n_29239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.202 0.0 33.23 0.163 ;
      END
   END n_29239

   PIN n_29241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.802 0.0 58.83 0.163 ;
      END
   END n_29241

   PIN n_29246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.442 0.0 59.47 0.163 ;
      END
   END n_29246

   PIN n_29249
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.482 0.0 58.51 0.163 ;
      END
   END n_29249

   PIN n_29264
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.402 0.0 60.43 0.163 ;
      END
   END n_29264

   PIN n_29280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.634 0.0 59.662 0.163 ;
      END
   END n_29280

   PIN n_29332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.01 0.0 57.038 0.163 ;
      END
   END n_29332

   PIN n_29350
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.162 0.0 58.19 0.163 ;
      END
   END n_29350

   PIN n_29362
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.754 0.0 32.782 0.163 ;
      END
   END n_29362

   PIN n_29371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.546 0.0 58.574 0.163 ;
      END
   END n_29371

   PIN n_29378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.394 0.0 57.422 0.163 ;
      END
   END n_29378

   PIN n_29461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.754 0.0 56.782 0.163 ;
      END
   END n_29461

   PIN n_29470
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.898 0.0 54.926 0.163 ;
      END
   END n_29470

   PIN n_29524
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.85 0.0 36.878 0.163 ;
      END
   END n_29524

   PIN n_29539
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.266 0.0 33.294 0.163 ;
      END
   END n_29539

   PIN n_29544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.586 0.0 57.614 0.163 ;
      END
   END n_29544

   PIN n_29549
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.834 0.0 54.862 0.163 ;
      END
   END n_29549

   PIN n_29562
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.074 0.0 33.102 0.163 ;
      END
   END n_29562

   PIN n_29593
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.562 0.0 32.59 0.163 ;
      END
   END n_29593

   PIN n_29594
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.818 0.0 24.846 0.163 ;
      END
   END n_29594

   PIN n_29595
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.498 0.0 32.526 0.163 ;
      END
   END n_29595

   PIN n_29611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.746 0.0 29.774 0.163 ;
      END
   END n_29611

   PIN n_29645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.626 0.0 24.654 0.163 ;
      END
   END n_29645

   PIN n_29649
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.746 0.0 29.774 0.163 ;
      END
   END n_29649

   PIN n_29753
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.538 0.0 63.566 0.163 ;
      END
   END n_29753

   PIN n_29756
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.01 0.0 33.038 0.163 ;
      END
   END n_29756

   PIN n_29817
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.69 0.0 40.718 0.163 ;
      END
   END n_29817

   PIN n_29840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.578 0.0 94.606 0.163 ;
      END
   END n_29840

   PIN n_29877
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.33 0.0 121.358 0.163 ;
      END
   END n_29877

   PIN n_29906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.658 0.0 108.686 0.163 ;
      END
   END n_29906

   PIN n_29918
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.274 0.0 36.302 0.163 ;
      END
   END n_29918

   PIN n_29943
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.242 0.0 56.27 0.163 ;
      END
   END n_29943

   PIN n_29949
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.314 0.0 107.342 0.163 ;
      END
   END n_29949

   PIN n_29998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 125.49 0.0 125.518 0.163 ;
      END
   END n_29998

   PIN n_30001
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.186 0.0 107.214 0.163 ;
      END
   END n_30001

   PIN n_30010
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.962 0.0 38.99 0.163 ;
      END
   END n_30010

   PIN n_30013
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.674 0.0 106.702 0.163 ;
      END
   END n_30013

   PIN n_30018
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.594 0.0 36.622 0.163 ;
      END
   END n_30018

   PIN n_30045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.746 0.0 109.774 0.163 ;
      END
   END n_30045

   PIN n_30049
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 129.266 0.0 129.294 0.163 ;
      END
   END n_30049

   PIN n_30051
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.586 0.0 121.614 0.163 ;
      END
   END n_30051

   PIN n_30107
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.834 0.0 118.862 0.163 ;
      END
   END n_30107

   PIN n_30111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.466 0.0 44.494 0.163 ;
      END
   END n_30111

   PIN n_30142
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.146 0.0 52.174 0.082 ;
      END
   END n_30142

   PIN n_30206
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.33 0.0 105.358 0.163 ;
      END
   END n_30206

   PIN n_30225
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.402 0.0 44.43 0.163 ;
      END
   END n_30225

   PIN n_30242
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.402 0.0 116.43 0.163 ;
      END
   END n_30242

   PIN n_30259
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.394 0.0 121.422 0.163 ;
      END
   END n_30259

   PIN n_30263
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.042 0.0 133.07 0.163 ;
      END
   END n_30263

   PIN n_30295
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.298 0.0 117.326 0.163 ;
      END
   END n_30295

   PIN n_30358
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.562 0.0 104.59 0.163 ;
      END
   END n_30358

   PIN n_30390
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.922 0.0 119.95 0.163 ;
      END
   END n_30390

   PIN n_30400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.714 0.0 113.742 0.163 ;
      END
   END n_30400

   PIN n_30406
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.65 0.0 113.678 0.163 ;
      END
   END n_30406

   PIN n_30418
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.394 0.0 121.422 0.163 ;
      END
   END n_30418

   PIN n_3045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.658 0.0 4.686 0.163 ;
      END
   END n_3045

   PIN n_30454
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.21 0.0 108.238 0.163 ;
      END
   END n_30454

   PIN n_30461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.546 0.0 106.574 0.163 ;
      END
   END n_30461

   PIN n_30527
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.026 0.0 119.054 0.163 ;
      END
   END n_30527

   PIN n_30528
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.25 0.0 115.278 0.163 ;
      END
   END n_30528

   PIN n_30544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.458 0.0 121.486 0.163 ;
      END
   END n_30544

   PIN n_30655
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.994 0.0 107.022 0.163 ;
      END
   END n_30655

   PIN n_30686
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 125.554 0.0 125.582 0.163 ;
      END
   END n_30686

   PIN n_30726
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.978 0.0 117.006 0.163 ;
      END
   END n_30726

   PIN n_30745
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 138.29 0.0 138.318 0.163 ;
      END
   END n_30745

   PIN n_30755
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.586 0.0 113.614 0.163 ;
      END
   END n_30755

   PIN n_30780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.458 0.0 121.486 0.163 ;
      END
   END n_30780

   PIN n_30792
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.65 0.0 121.678 0.163 ;
      END
   END n_30792

   PIN n_30818
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.562 0.0 40.59 0.082 ;
      END
   END n_30818

   PIN n_30835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.106 0.0 133.134 0.163 ;
      END
   END n_30835

   PIN n_30917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.298 0.0 109.326 0.163 ;
      END
   END n_30917

   PIN n_30997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.306 0.0 120.334 0.163 ;
      END
   END n_30997

   PIN n_31021
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.714 0.0 121.742 0.163 ;
      END
   END n_31021

   PIN n_31023
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.122 0.0 115.15 0.163 ;
      END
   END n_31023

   PIN n_31039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.49 0.0 125.518 0.163 ;
      END
   END n_31039

   PIN n_31077
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.482 0.0 106.51 0.163 ;
      END
   END n_31077

   PIN n_31091
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.194 0.0 110.222 0.163 ;
      END
   END n_31091

   PIN n_31095
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.418 0.0 114.446 0.163 ;
      END
   END n_31095

   PIN n_31106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.978 0.0 45.006 0.163 ;
      END
   END n_31106

   PIN n_31114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.434 0.0 40.462 0.163 ;
      END
   END n_31114

   PIN n_31122
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 125.618 0.0 125.646 0.163 ;
      END
   END n_31122

   PIN n_31130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 46.77 0.0 46.798 0.163 ;
      END
   END n_31130

   PIN n_31132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.098 0.0 114.126 0.163 ;
      END
   END n_31132

   PIN n_31146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.658 0.0 108.686 0.163 ;
      END
   END n_31146

   PIN n_31149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.554 0.0 109.582 0.163 ;
      END
   END n_31149

   PIN n_31165
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.658 0.0 44.686 0.163 ;
      END
   END n_31165

   PIN n_31179
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.754 0.0 40.782 0.163 ;
      END
   END n_31179

   PIN n_31222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.266 0.0 129.294 0.163 ;
      END
   END n_31222

   PIN n_31280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.682 0.0 109.71 0.163 ;
      END
   END n_31280

   PIN n_31288
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.73 0.0 55.758 0.163 ;
      END
   END n_31288

   PIN n_31304
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.722 0.0 108.75 0.163 ;
      END
   END n_31304

   PIN n_31306
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.106 0.0 109.134 0.163 ;
      END
   END n_31306

   PIN n_31333
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 46.642 0.0 46.67 0.163 ;
      END
   END n_31333

   PIN n_31342
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.29 0.0 42.318 0.163 ;
      END
   END n_31342

   PIN n_31345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.434 0.0 40.462 0.163 ;
      END
   END n_31345

   PIN n_3136
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.402 0.163 20.43 ;
      END
   END n_3136

   PIN n_31381
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.226 0.0 42.254 0.163 ;
      END
   END n_31381

   PIN n_31430
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.306 0.0 48.334 0.163 ;
      END
   END n_31430

   PIN n_31463
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.69 0.0 40.718 0.163 ;
      END
   END n_31463

   PIN n_31464
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.266 0.0 105.294 0.163 ;
      END
   END n_31464

   PIN n_31479
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.722 0.0 44.75 0.163 ;
      END
   END n_31479

   PIN n_31497
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.794 0.0 103.822 0.163 ;
      END
   END n_31497

   PIN n_31510
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.33 0.0 113.358 0.163 ;
      END
   END n_31510

   PIN n_31514
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.066 0.0 46.094 0.163 ;
      END
   END n_31514

   PIN n_31533
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.978 0.0 37.006 0.163 ;
      END
   END n_31533

   PIN n_31543
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.93 0.0 114.958 0.163 ;
      END
   END n_31543

   PIN n_31544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.866 0.0 114.894 0.163 ;
      END
   END n_31544

   PIN n_31547
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.842 0.0 113.87 0.163 ;
      END
   END n_31547

   PIN n_31552
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.066 0.0 110.094 0.163 ;
      END
   END n_31552

   PIN n_31587
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.37 0.0 40.398 0.163 ;
      END
   END n_31587

   PIN n_31609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.306 0.0 40.334 0.163 ;
      END
   END n_31609

   PIN n_31644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.69 0.0 48.718 0.163 ;
      END
   END n_31644

   PIN n_3165
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.954 0.163 3.982 ;
      END
   END n_3165

   PIN n_31657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.514 0.0 110.542 0.163 ;
      END
   END n_31657

   PIN n_31659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.658 0.0 44.686 0.163 ;
      END
   END n_31659

   PIN n_31667
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.242 0.0 40.27 0.163 ;
      END
   END n_31667

   PIN n_31668
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.466 0.0 44.494 0.163 ;
      END
   END n_31668

   PIN n_31669
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.402 0.0 44.43 0.163 ;
      END
   END n_31669

   PIN n_31684
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.45 0.0 110.478 0.163 ;
      END
   END n_31684

   PIN n_31685
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.802 0.0 74.83 0.163 ;
      END
   END n_31685

   PIN n_31701
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.802 0.0 98.83 0.163 ;
      END
   END n_31701

   PIN n_31716
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.21 0.0 100.238 0.163 ;
      END
   END n_31716

   PIN n_31733
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.53 0.0 44.558 0.163 ;
      END
   END n_31733

   PIN n_31742
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.682 0.0 85.71 0.163 ;
      END
   END n_31742

   PIN n_31745
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.25 0.0 83.278 0.163 ;
      END
   END n_31745

   PIN n_31829
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.442 0.0 51.47 0.163 ;
      END
   END n_31829

   PIN n_31855
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.362 0.0 69.39 0.163 ;
      END
   END n_31855

   PIN n_31857
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.282 0.0 71.31 0.163 ;
      END
   END n_31857

   PIN n_3189
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.37 0.163 8.398 ;
      END
   END n_3189

   PIN n_31896
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.018 0.0 52.046 0.163 ;
      END
   END n_31896

   PIN n_31898
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 68.466 0.0 68.494 0.163 ;
      END
   END n_31898

   PIN n_31911
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.306 0.0 64.334 0.163 ;
      END
   END n_31911

   PIN n_32023
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.89 0.0 99.918 0.163 ;
      END
   END n_32023

   PIN n_32055
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.282 0.0 79.31 0.163 ;
      END
   END n_32055

   PIN n_32071
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.354 0.0 66.382 0.163 ;
      END
   END n_32071

   PIN n_32181
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.154 0.0 55.182 0.163 ;
      END
   END n_32181

   PIN n_32200
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.338 0.0 68.366 0.163 ;
      END
   END n_32200

   PIN n_32218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.058 0.0 83.086 0.163 ;
      END
   END n_32218

   PIN n_32268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.89 0.0 67.918 0.163 ;
      END
   END n_32268

   PIN n_32272
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.986 0.0 64.014 0.163 ;
      END
   END n_32272

   PIN n_32333
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.01 0.0 65.038 0.163 ;
      END
   END n_32333

   PIN n_32511
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.042 0.0 69.07 0.163 ;
      END
   END n_32511

   PIN n_32526
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.418 0.0 42.446 0.163 ;
      END
   END n_32526

   PIN n_32586
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.418 0.0 66.446 0.163 ;
      END
   END n_32586

   PIN n_32608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.506 0.0 43.534 0.163 ;
      END
   END n_32608

   PIN n_32620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.882 0.0 64.91 0.163 ;
      END
   END n_32620

   PIN n_32650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.73 0.0 71.758 0.163 ;
      END
   END n_32650

   PIN n_32654
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.874 0.0 69.902 0.163 ;
      END
   END n_32654

   PIN n_32662
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.946 0.0 64.974 0.163 ;
      END
   END n_32662

   PIN n_32677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.946 0.0 64.974 0.163 ;
      END
   END n_32677

   PIN n_32678
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.058 0.0 83.086 0.163 ;
      END
   END n_32678

   PIN n_32695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.922 0.0 71.95 0.163 ;
      END
   END n_32695

   PIN n_32766
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.986 0.0 72.014 0.163 ;
      END
   END n_32766

   PIN n_32777
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.434 0.0 48.462 0.163 ;
      END
   END n_32777

   PIN n_32803
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.618 0.0 69.646 0.163 ;
      END
   END n_32803

   PIN n_32804
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 72.498 0.0 72.526 0.163 ;
      END
   END n_32804

   PIN n_32807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.09 0.0 71.118 0.163 ;
      END
   END n_32807

   PIN n_32810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.858 0.0 63.886 0.163 ;
      END
   END n_32810

   PIN n_32811
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.754 0.0 48.782 0.163 ;
      END
   END n_32811

   PIN n_32828
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.354 0.0 66.382 0.163 ;
      END
   END n_32828

   PIN n_32865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.29 0.0 66.318 0.163 ;
      END
   END n_32865

   PIN n_32866
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.938 0.0 101.966 0.082 ;
      END
   END n_32866

   PIN n_32927
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.162 0.0 66.19 0.163 ;
      END
   END n_32927

   PIN n_32952
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.914 0.0 68.942 0.163 ;
      END
   END n_32952

   PIN n_32970
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.282 0.0 63.31 0.163 ;
      END
   END n_32970

   PIN n_32976
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.346 0.0 63.374 0.163 ;
      END
   END n_32976

   PIN n_33002
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.378 0.0 75.406 0.163 ;
      END
   END n_33002

   PIN n_33019
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.306 0.0 64.334 0.163 ;
      END
   END n_33019

   PIN n_33073
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.194 0.0 70.222 0.163 ;
      END
   END n_33073

   PIN n_33080
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.69 0.0 72.718 0.163 ;
      END
   END n_33080

   PIN n_33098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.258 0.0 70.286 0.163 ;
      END
   END n_33098

   PIN n_33134
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.866 0.0 66.894 0.163 ;
      END
   END n_33134

   PIN n_33154
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.41 0.0 63.438 0.163 ;
      END
   END n_33154

   PIN n_33172
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.69 0.0 48.718 0.163 ;
      END
   END n_33172

   PIN n_33210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.386 0.0 70.414 0.163 ;
      END
   END n_33210

   PIN n_33229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.57 0.0 67.598 0.163 ;
      END
   END n_33229

   PIN n_33295
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.026 0.0 71.054 0.163 ;
      END
   END n_33295

   PIN n_33371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.738 0.0 66.766 0.163 ;
      END
   END n_33371

   PIN n_33389
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.626 0.0 48.654 0.163 ;
      END
   END n_33389

   PIN n_33406
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.354 0.0 42.382 0.163 ;
      END
   END n_33406

   PIN n_33437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.698 0.0 43.726 0.163 ;
      END
   END n_33437

   PIN n_33472
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.762 0.0 43.79 0.163 ;
      END
   END n_33472

   PIN n_33499
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.866 0.0 42.894 0.163 ;
      END
   END n_33499

   PIN n_3351
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.098 0.163 10.126 ;
      END
   END n_3351

   PIN n_33543
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.666 0.0 63.694 0.163 ;
      END
   END n_33543

   PIN n_33601
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.922 0.0 39.95 0.163 ;
      END
   END n_33601

   PIN n_33602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.594 0.0 44.622 0.163 ;
      END
   END n_33602

   PIN n_33603
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.594 0.0 44.622 0.163 ;
      END
   END n_33603

   PIN n_33604
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.53 0.0 44.558 0.163 ;
      END
   END n_33604

   PIN n_33627
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 80.626 0.0 80.654 0.163 ;
      END
   END n_33627

   PIN n_33638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.474 0.0 63.502 0.163 ;
      END
   END n_33638

   PIN n_33667
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.282 0.0 63.31 0.163 ;
      END
   END n_33667

   PIN n_33701
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.218 0.0 63.246 0.163 ;
      END
   END n_33701

   PIN n_33735
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.274 0.0 52.302 0.163 ;
      END
   END n_33735

   PIN n_33977
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.026 0.0 87.054 0.163 ;
      END
   END n_33977

   PIN n_34040
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.402 0.0 92.43 0.163 ;
      END
   END n_34040

   PIN n_34127
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.378 0.0 91.406 0.163 ;
      END
   END n_34127

   PIN n_34204
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.354 0.0 90.382 0.163 ;
      END
   END n_34204

   PIN n_34217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.09 0.0 95.118 0.163 ;
      END
   END n_34217

   PIN n_34298
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.25 0.0 83.278 0.163 ;
      END
   END n_34298

   PIN n_34312
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.65 0.0 89.678 0.163 ;
      END
   END n_34312

   PIN n_34315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.186 0.0 91.214 0.163 ;
      END
   END n_34315

   PIN n_34369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.218 0.0 87.246 0.163 ;
      END
   END n_34369

   PIN n_34418
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.746 0.0 93.774 0.163 ;
      END
   END n_34418

   PIN n_34420
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.97 0.0 89.998 0.163 ;
      END
   END n_34420

   PIN n_34475
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.082 0.0 92.11 0.163 ;
      END
   END n_34475

   PIN n_34501
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.77 0.0 86.798 0.163 ;
      END
   END n_34501

   PIN n_34505
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.29 0.0 90.318 0.082 ;
      END
   END n_34505

   PIN n_3452
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.482 0.163 10.51 ;
      END
   END n_3452

   PIN n_34605
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.546 0.0 90.574 0.163 ;
      END
   END n_34605

   PIN n_34738
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.642 0.0 86.67 0.163 ;
      END
   END n_34738

   PIN n_34794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.57 0.0 91.598 0.163 ;
      END
   END n_34794

   PIN n_34839
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.218 0.0 95.246 0.163 ;
      END
   END n_34839

   PIN n_34903
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.578 0.0 94.606 0.163 ;
      END
   END n_34903

   PIN n_34918
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.026 0.0 95.054 0.163 ;
      END
   END n_34918

   PIN n_34999
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.146 0.0 92.174 0.163 ;
      END
   END n_34999

   PIN n_35106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.898 0.0 94.926 0.163 ;
      END
   END n_35106

   PIN n_35141
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.93 0.0 90.958 0.163 ;
      END
   END n_35141

   PIN n_35319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.946 0.0 88.974 0.163 ;
      END
   END n_35319

   PIN n_3533
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.05 0.163 24.078 ;
      END
   END n_3533

   PIN n_35567
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.794 0.0 95.822 0.163 ;
      END
   END n_35567

   PIN n_3607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.466 0.163 20.494 ;
      END
   END n_3607

   PIN n_3623
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.018 0.163 4.046 ;
      END
   END n_3623

   PIN n_3863
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.314 0.163 3.342 ;
      END
   END n_3863

   PIN n_3903
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.034 0.0 2.062 0.163 ;
      END
   END n_3903

   PIN n_3909
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.738 0.0 2.766 0.163 ;
      END
   END n_3909

   PIN n_3935
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.25 0.163 3.278 ;
      END
   END n_3935

   PIN n_4062
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.138 0.0 1.166 0.163 ;
      END
   END n_4062

   PIN n_4064
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.53 0.163 20.558 ;
      END
   END n_4064

   PIN n_4068
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.306 0.163 8.334 ;
      END
   END n_4068

   PIN n_4079
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.186 0.163 3.214 ;
      END
   END n_4079

   PIN n_4088
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.082 0.0 4.11 0.163 ;
      END
   END n_4088

   PIN n_4104
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.578 0.163 6.606 ;
      END
   END n_4104

   PIN n_4105
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.202 0.0 9.23 0.163 ;
      END
   END n_4105

   PIN n_4118
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.546 0.163 10.574 ;
      END
   END n_4118

   PIN n_4122
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.906 0.0 9.934 0.163 ;
      END
   END n_4122

   PIN n_4131
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.13 0.0 6.158 0.163 ;
      END
   END n_4131

   PIN n_4201
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.594 0.163 20.622 ;
      END
   END n_4201

   PIN n_4204
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.842 0.0 9.87 0.163 ;
      END
   END n_4204

   PIN n_4294
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.074 0.0 1.102 0.163 ;
      END
   END n_4294

   PIN n_4490
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.354 0.0 2.382 0.163 ;
      END
   END n_4490

   PIN n_4494
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.61 0.0 2.638 0.163 ;
      END
   END n_4494

   PIN n_4561
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.37 0.0 0.398 0.163 ;
      END
   END n_4561

   PIN n_4708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.994 0.0 11.022 0.163 ;
      END
   END n_4708

   PIN n_4799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.634 0.163 3.662 ;
      END
   END n_4799

   PIN n_4811
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.65 0.0 1.678 0.163 ;
      END
   END n_4811

   PIN n_4882
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.962 0.163 6.99 ;
      END
   END n_4882

   PIN n_4923
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.866 0.0 2.894 0.163 ;
      END
   END n_4923

   PIN n_4958
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.178 0.0 8.206 0.163 ;
      END
   END n_4958

   PIN n_4961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.986 0.163 16.014 ;
      END
   END n_4961

   PIN n_5049
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.05 0.163 16.078 ;
      END
   END n_5049

   PIN n_5069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.61 0.0 10.638 0.163 ;
      END
   END n_5069

   PIN n_5268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.474 0.0 7.502 0.163 ;
      END
   END n_5268

   PIN n_5314
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.97 0.0 9.998 0.163 ;
      END
   END n_5314

   PIN n_5323
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.234 0.0 13.262 0.163 ;
      END
   END n_5323

   PIN n_5363
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.794 0.0 7.822 0.163 ;
      END
   END n_5363

   PIN n_5372
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.114 0.163 24.142 ;
      END
   END n_5372

   PIN n_5437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.018 0.0 12.046 0.163 ;
      END
   END n_5437

   PIN n_5482
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.426 0.0 13.454 0.163 ;
      END
   END n_5482

   PIN n_5571
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.026 0.0 15.054 0.163 ;
      END
   END n_5571

   PIN n_5574
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.306 0.163 24.334 ;
      END
   END n_5574

   PIN n_5581
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.082 0.163 12.11 ;
      END
   END n_5581

   PIN n_5643
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.402 0.0 12.43 0.163 ;
      END
   END n_5643

   PIN n_59574
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.226 0.163 10.254 ;
      END
   END n_59574

   PIN n_6096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.994 0.0 19.022 0.163 ;
      END
   END n_6096

   PIN n_61534
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.466 0.163 4.494 ;
      END
   END n_61534

   PIN n_61611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.754 0.0 0.782 0.163 ;
      END
   END n_61611

   PIN n_6257
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.53 0.0 12.558 0.163 ;
      END
   END n_6257

   PIN n_63161
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.882 0.163 8.91 ;
      END
   END n_63161

   PIN n_63230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.106 94.557 37.134 94.72 ;
      END
   END n_63230

   PIN n_63234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.906 0.163 9.934 ;
      END
   END n_63234

   PIN n_63421
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.122 0.163 11.15 ;
      END
   END n_63421

   PIN n_63508
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.506 0.0 3.534 0.163 ;
      END
   END n_63508

   PIN n_63603
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.49 0.0 21.518 0.163 ;
      END
   END n_63603

   PIN n_63622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.93 0.163 58.958 ;
      END
   END n_63622

   PIN n_63690
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 32.626 0.163 32.654 ;
      END
   END n_63690

   PIN n_63695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.21 0.163 28.238 ;
      END
   END n_63695

   PIN n_63776
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.738 0.163 58.766 ;
      END
   END n_63776

   PIN n_63794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.914 0.0 20.942 0.163 ;
      END
   END n_63794

   PIN n_63840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.538 0.0 23.566 0.163 ;
      END
   END n_63840

   PIN n_63851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.834 0.0 22.862 0.163 ;
      END
   END n_63851

   PIN n_63858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.09 0.0 23.118 0.082 ;
      END
   END n_63858

   PIN n_63883
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.602 0.0 23.63 0.163 ;
      END
   END n_63883

   PIN n_63885
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.05 0.0 24.078 0.163 ;
      END
   END n_63885

   PIN n_63886
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.282 0.0 23.31 0.163 ;
      END
   END n_63886

   PIN n_63972
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.85 0.0 20.878 0.163 ;
      END
   END n_63972

   PIN n_64022
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.578 0.0 22.606 0.163 ;
      END
   END n_64022

   PIN n_64028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.346 0.163 47.374 ;
      END
   END n_64028

   PIN n_64034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.17 0.0 5.198 0.163 ;
      END
   END n_64034

   PIN n_64049
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.81 0.0 21.838 0.163 ;
      END
   END n_64049

   PIN n_64091
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 28.146 0.163 28.174 ;
      END
   END n_64091

   PIN n_64119
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 32.754 0.082 32.782 ;
      END
   END n_64119

   PIN n_64138
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.658 0.0 20.686 0.163 ;
      END
   END n_64138

   PIN n_64153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.922 0.163 31.95 ;
      END
   END n_64153

   PIN n_64188
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.866 0.163 58.894 ;
      END
   END n_64188

   PIN n_64189
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.802 0.163 58.83 ;
      END
   END n_64189

   PIN n_64248
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.09 0.0 23.118 0.163 ;
      END
   END n_64248

   PIN n_64308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 28.21 0.163 28.238 ;
      END
   END n_64308

   PIN n_64341
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.674 0.163 58.702 ;
      END
   END n_64341

   PIN n_64388
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.026 0.0 23.054 0.163 ;
      END
   END n_64388

   PIN n_64414
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.858 0.163 31.886 ;
      END
   END n_64414

   PIN n_64439
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.986 0.0 24.014 0.163 ;
      END
   END n_64439

   PIN n_64590
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.554 0.0 21.582 0.163 ;
      END
   END n_64590

   PIN n_64618
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.946 0.0 24.974 0.163 ;
      END
   END n_64618

   PIN n_64713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.882 0.0 24.91 0.163 ;
      END
   END n_64713

   PIN n_64732
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.514 0.0 22.542 0.163 ;
      END
   END n_64732

   PIN n_64733
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.818 0.0 24.846 0.163 ;
      END
   END n_64733

   PIN n_64736
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.682 0.0 21.71 0.163 ;
      END
   END n_64736

   PIN n_64749
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.962 0.0 22.99 0.163 ;
      END
   END n_64749

   PIN n_64824
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.978 0.0 21.006 0.163 ;
      END
   END n_64824

   PIN n_64842
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.626 0.0 24.654 0.163 ;
      END
   END n_64842

   PIN n_64909
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.85 0.0 20.878 0.163 ;
      END
   END n_64909

   PIN n_64922
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.082 0.0 20.11 0.163 ;
      END
   END n_64922

   PIN n_64923
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.786 0.0 20.814 0.163 ;
      END
   END n_64923

   PIN n_64962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.514 0.163 62.542 ;
      END
   END n_64962

   PIN n_65028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.81 0.0 29.838 0.163 ;
      END
   END n_65028

   PIN n_6503
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.618 0.0 61.646 0.163 ;
      END
   END n_6503

   PIN n_65155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.466 0.0 20.494 0.163 ;
      END
   END n_65155

   PIN n_65446
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.642 0.0 6.67 0.163 ;
      END
   END n_65446

   PIN n_65451
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.77 0.0 6.798 0.163 ;
      END
   END n_65451

   PIN n_65473
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.73 0.163 39.758 ;
      END
   END n_65473

   PIN n_65475
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.826 0.0 27.854 0.163 ;
      END
   END n_65475

   PIN n_65507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.234 0.163 13.262 ;
      END
   END n_65507

   PIN n_65527
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.378 0.082 11.406 ;
      END
   END n_65527

   PIN n_65552
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.162 0.163 10.19 ;
      END
   END n_65552

   PIN n_65560
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.21 0.0 12.238 0.163 ;
      END
   END n_65560

   PIN n_65578
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.154 0.0 15.182 0.163 ;
      END
   END n_65578

   PIN n_65583
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.49 0.163 13.518 ;
      END
   END n_65583

   PIN n_65610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.274 0.163 12.302 ;
      END
   END n_65610

   PIN n_65621
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.81 0.163 13.838 ;
      END
   END n_65621

   PIN n_65671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.378 0.0 27.406 0.163 ;
      END
   END n_65671

   PIN n_65702
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.218 0.0 15.246 0.163 ;
      END
   END n_65702

   PIN n_65747
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.282 0.0 15.31 0.163 ;
      END
   END n_65747

   PIN n_65752
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.354 0.0 26.382 0.163 ;
      END
   END n_65752

   PIN n_65753
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.402 0.163 4.43 ;
      END
   END n_65753

   PIN n_65810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.466 0.163 12.494 ;
      END
   END n_65810

   PIN n_65890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.114 0.163 16.142 ;
      END
   END n_65890

   PIN n_65897
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.954 0.163 11.982 ;
      END
   END n_65897

   PIN n_65923
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.034 0.0 26.062 0.163 ;
      END
   END n_65923

   PIN n_65941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.29 0.163 10.318 ;
      END
   END n_65941

   PIN n_65953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.338 0.163 12.366 ;
      END
   END n_65953

   PIN n_65962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.482 0.0 26.51 0.163 ;
      END
   END n_65962

   PIN n_65965
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.61 0.0 26.638 0.163 ;
      END
   END n_65965

   PIN n_65979
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.178 0.163 16.206 ;
      END
   END n_65979

   PIN n_66001
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.898 0.0 14.926 0.163 ;
      END
   END n_66001

   PIN n_66004
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.194 0.0 14.222 0.163 ;
      END
   END n_66004

   PIN n_66070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.442 0.0 27.47 0.163 ;
      END
   END n_66070

   PIN n_66106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.146 0.163 12.174 ;
      END
   END n_66106

   PIN n_66122
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.114 0.0 16.142 0.163 ;
      END
   END n_66122

   PIN n_66130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.434 0.163 16.462 ;
      END
   END n_66130

   PIN n_66184
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.842 0.0 25.87 0.163 ;
      END
   END n_66184

   PIN n_66209
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.97 0.0 25.998 0.163 ;
      END
   END n_66209

   PIN n_66223
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.162 0.0 26.19 0.163 ;
      END
   END n_66223

   PIN n_66292
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.058 0.0 27.086 0.163 ;
      END
   END n_66292

   PIN n_66319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.946 94.557 40.974 94.72 ;
      END
   END n_66319

   PIN n_66357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.386 0.0 14.414 0.163 ;
      END
   END n_66357

   PIN n_66374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.458 0.0 25.486 0.082 ;
      END
   END n_66374

   PIN n_66380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.954 0.163 3.982 ;
      END
   END n_66380

   PIN n_66389
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 0.0 25.614 0.163 ;
      END
   END n_66389

   PIN n_66417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.178 0.163 16.206 ;
      END
   END n_66417

   PIN n_66438
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.89 0.163 3.918 ;
      END
   END n_66438

   PIN n_66469
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.906 0.0 25.934 0.163 ;
      END
   END n_66469

   PIN n_66475
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.554 0.0 13.582 0.163 ;
      END
   END n_66475

   PIN n_66487
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.25 0.163 11.278 ;
      END
   END n_66487

   PIN n_66506
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.106 0.0 29.134 0.163 ;
      END
   END n_66506

   PIN n_66569
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.978 0.0 13.006 0.163 ;
      END
   END n_66569

   PIN n_66584
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.938 0.0 13.966 0.163 ;
      END
   END n_66584

   PIN n_66589
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.426 0.0 13.454 0.163 ;
      END
   END n_66589

   PIN n_66623
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.89 0.163 11.918 ;
      END
   END n_66623

   PIN n_66630
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.826 0.163 11.854 ;
      END
   END n_66630

   PIN n_66656
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.794 0.163 31.822 ;
      END
   END n_66656

   PIN n_66678
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.514 0.0 14.542 0.163 ;
      END
   END n_66678

   PIN n_66807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.242 0.0 0.27 0.163 ;
      END
   END n_66807

   PIN n_66822
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.698 0.163 35.726 ;
      END
   END n_66822

   PIN n_66873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.762 0.163 11.79 ;
      END
   END n_66873

   PIN n_67053
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.418 0.163 10.446 ;
      END
   END n_67053

   PIN n_67065
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.882 94.557 40.91 94.72 ;
      END
   END n_67065

   PIN n_67119
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.698 0.163 11.726 ;
      END
   END n_67119

   PIN n_67131
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.034 94.557 18.062 94.72 ;
      END
   END n_67131

   PIN n_67150
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.666 0.163 39.694 ;
      END
   END n_67150

   PIN n_67203
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.314 0.163 3.342 ;
      END
   END n_67203

   PIN n_67231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.602 0.163 39.63 ;
      END
   END n_67231

   PIN n_67232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.538 0.163 39.566 ;
      END
   END n_67232

   PIN n_67245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.226 94.557 42.254 94.72 ;
      END
   END n_67245

   PIN n_67246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.754 94.557 40.782 94.72 ;
      END
   END n_67246

   PIN n_67247
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.106 94.557 37.134 94.72 ;
      END
   END n_67247

   PIN n_67326
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.906 94.557 17.934 94.72 ;
      END
   END n_67326

   PIN n_67480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.546 0.0 18.574 0.163 ;
      END
   END n_67480

   PIN n_67630
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.33 0.0 17.358 0.082 ;
      END
   END n_67630

   PIN n_67644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.522 0.0 17.55 0.163 ;
      END
   END n_67644

   PIN n_67654
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.538 0.0 15.566 0.163 ;
      END
   END n_67654

   PIN n_67771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.61 0.0 18.638 0.163 ;
      END
   END n_67771

   PIN n_67793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.906 0.0 17.934 0.163 ;
      END
   END n_67793

   PIN n_67946
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.69 0.0 16.718 0.163 ;
      END
   END n_67946

   PIN n_67996
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.562 0.0 40.59 0.163 ;
      END
   END n_67996

   PIN n_68009
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.202 0.0 17.23 0.163 ;
      END
   END n_68009

   PIN n_68020
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.146 0.163 28.174 ;
      END
   END n_68020

   PIN n_68045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.354 0.0 18.382 0.163 ;
      END
   END n_68045

   PIN n_68057
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.082 0.163 28.11 ;
      END
   END n_68057

   PIN n_68205
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.474 0.0 15.502 0.163 ;
      END
   END n_68205

   PIN n_68264
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.042 0.0 29.07 0.163 ;
      END
   END n_68264

   PIN n_68269
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.626 0.0 16.654 0.163 ;
      END
   END n_68269

   PIN n_68283
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.33 0.0 17.358 0.163 ;
      END
   END n_68283

   PIN n_68286
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.602 0.0 15.63 0.163 ;
      END
   END n_68286

   PIN n_68349
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.074 0.0 25.102 0.163 ;
      END
   END n_68349

   PIN n_68352
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.97 0.0 17.998 0.163 ;
      END
   END n_68352

   PIN n_68366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.458 0.0 17.486 0.163 ;
      END
   END n_68366

   PIN n_68377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.122 0.0 19.15 0.163 ;
      END
   END n_68377

   PIN n_68515
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.09 0.0 15.118 0.163 ;
      END
   END n_68515

   PIN n_68805
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.138 0.0 17.166 0.163 ;
      END
   END n_68805

   PIN n_69023
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.242 0.163 24.27 ;
      END
   END n_69023

   PIN n_69052
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.178 0.163 24.206 ;
      END
   END n_69052

   PIN n_69101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.018 0.163 28.046 ;
      END
   END n_69101

   PIN n_69155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.858 0.163 15.886 ;
      END
   END n_69155

   PIN n_69285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.274 0.163 12.302 ;
      END
   END n_69285

   PIN n_6944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.49 0.0 29.518 0.163 ;
      END
   END n_6944

   PIN n_69515
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.65 0.0 17.678 0.163 ;
      END
   END n_69515

   PIN n_69551
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.37 0.163 16.398 ;
      END
   END n_69551

   PIN n_69624
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.106 0.0 21.134 0.163 ;
      END
   END n_69624

   PIN n_69650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.698 0.0 11.726 0.163 ;
      END
   END n_69650

   PIN n_69668
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.378 0.0 11.406 0.082 ;
      END
   END n_69668

   PIN n_69677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.098 0.0 98.126 0.163 ;
      END
   END n_69677

   PIN n_69697
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.826 0.0 11.854 0.163 ;
      END
   END n_69697

   PIN n_69698
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.194 0.0 22.222 0.163 ;
      END
   END n_69698

   PIN n_69751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.554 0.0 29.582 0.163 ;
      END
   END n_69751

   PIN n_69798
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.162 0.0 106.19 0.163 ;
      END
   END n_69798

   PIN n_69817
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.29 0.0 18.318 0.163 ;
      END
   END n_69817

   PIN n_69828
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.13 0.0 22.158 0.163 ;
      END
   END n_69828

   PIN n_69839
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.17 0.0 21.198 0.163 ;
      END
   END n_69839

   PIN n_70031
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.034 0.0 98.062 0.163 ;
      END
   END n_70031

   PIN n_70168
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.002 0.0 110.03 0.163 ;
      END
   END n_70168

   PIN n_70237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.25 0.0 11.278 0.163 ;
      END
   END n_70237

   PIN n_70400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.97 0.0 105.998 0.163 ;
      END
   END n_70400

   PIN n_70401
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.29 0.0 106.318 0.163 ;
      END
   END n_70401

   PIN n_70488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.226 0.0 106.254 0.163 ;
      END
   END n_70488

   PIN n_70529
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.098 0.0 98.126 0.082 ;
      END
   END n_70529

   PIN n_70631
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.13 0.0 94.158 0.163 ;
      END
   END n_70631

   PIN n_70788
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.386 0.0 102.414 0.163 ;
      END
   END n_70788

   PIN n_7085
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.338 0.163 4.366 ;
      END
   END n_7085

   PIN n_70959
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.018 0.0 100.046 0.082 ;
      END
   END n_70959

   PIN n_70968
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.322 0.0 102.35 0.163 ;
      END
   END n_70968

   PIN n_70996
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.61 0.0 106.638 0.163 ;
      END
   END n_70996

   PIN n_71009
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.29 0.0 98.318 0.163 ;
      END
   END n_71009

   PIN n_71083
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.322 0.0 102.35 0.163 ;
      END
   END n_71083

   PIN n_71095
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.226 0.0 98.254 0.163 ;
      END
   END n_71095

   PIN n_71105
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.258 0.0 102.286 0.163 ;
      END
   END n_71105

   PIN n_71108
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.546 0.0 106.574 0.163 ;
      END
   END n_71108

   PIN n_71151
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.258 0.0 102.286 0.163 ;
      END
   END n_71151

   PIN n_71192
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.194 0.0 102.222 0.163 ;
      END
   END n_71192

   PIN n_7212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.946 0.0 48.974 0.163 ;
      END
   END n_7212

   PIN n_753
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.21 0.163 12.238 ;
      END
   END n_753

   PIN n_75355
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.546 0.0 10.574 0.163 ;
      END
   END n_75355

   PIN n_75387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.498 0.0 24.526 0.082 ;
      END
   END n_75387

   PIN n_75701
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.298 0.0 13.326 0.163 ;
      END
   END n_75701

   PIN n_75702
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.362 0.0 13.39 0.163 ;
      END
   END n_75702

   PIN n_75837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.586 0.0 17.614 0.163 ;
      END
   END n_75837

   PIN n_75950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.93 0.0 10.958 0.082 ;
      END
   END n_75950

   PIN n_75954
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.146 0.163 12.174 ;
      END
   END n_75954

   PIN n_76207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 17.01 0.163 17.038 ;
      END
   END n_76207

   PIN n_76269
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.69 0.0 24.718 0.163 ;
      END
   END n_76269

   PIN n_76439
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.754 0.0 8.782 0.163 ;
      END
   END n_76439

   PIN n_76451
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.122 0.0 11.15 0.163 ;
      END
   END n_76451

   PIN n_76463
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.466 0.0 4.494 0.163 ;
      END
   END n_76463

   PIN n_76471
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.546 0.0 10.574 0.163 ;
      END
   END n_76471

   PIN n_76474
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.114 0.163 16.142 ;
      END
   END n_76474

   PIN n_76570
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.482 0.0 10.51 0.163 ;
      END
   END n_76570

   PIN n_76637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.034 0.0 10.062 0.163 ;
      END
   END n_76637

   PIN n_76642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 17.074 0.163 17.102 ;
      END
   END n_76642

   PIN n_76809
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.058 0.0 11.086 0.163 ;
      END
   END n_76809

   PIN n_76821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.786 0.163 20.814 ;
      END
   END n_76821

   PIN n_77030
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 17.138 0.163 17.166 ;
      END
   END n_77030

   PIN n_77046
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.818 0.0 8.846 0.163 ;
      END
   END n_77046

   PIN n_77228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.658 0.163 20.686 ;
      END
   END n_77228

   PIN n_77801
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.722 0.163 20.75 ;
      END
   END n_77801

   PIN n_78115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.81 0.0 13.838 0.163 ;
      END
   END n_78115

   PIN n_7851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.746 0.0 5.774 0.163 ;
      END
   END n_7851

   PIN n_7898
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.818 0.0 0.846 0.163 ;
      END
   END n_7898

   PIN n_90978
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.818 0.0 120.846 0.163 ;
      END
   END n_90978

   PIN n_95123
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.202 0.0 81.23 0.163 ;
      END
   END n_95123

   PIN n_9943
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.266 0.0 9.294 0.163 ;
      END
   END n_9943

   PIN stage1_out_3187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.122 0.0 83.15 0.163 ;
      END
   END stage1_out_3187

   PIN stage1_out_3201
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.754 0.0 48.782 0.163 ;
      END
   END stage1_out_3201

   PIN stage1_out_3213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.866 0.0 18.894 0.163 ;
      END
   END stage1_out_3213

   PIN u0_IP_64__1299
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.682 94.557 21.71 94.72 ;
      END
   END u0_IP_64__1299

   PIN u0_L4_29_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.122 0.163 11.15 ;
      END
   END u0_L4_29_

   PIN u0_L5_30_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.986 0.163 24.014 ;
      END
   END u0_L5_30_

   PIN u0_L6_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.922 0.163 7.95 ;
      END
   END u0_L6_10_

   PIN u0_L6_21_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.362 0.0 29.39 0.163 ;
      END
   END u0_L6_21_

   PIN u0_L6_29_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.786 0.0 44.814 0.163 ;
      END
   END u0_L6_29_

   PIN u0_L7_20_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.642 0.0 94.67 0.163 ;
      END
   END u0_L7_20_

   PIN u0_L7_28_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.882 0.0 48.91 0.163 ;
      END
   END u0_L7_28_

   PIN u0_L8_20_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.706 0.0 94.734 0.163 ;
      END
   END u0_L8_20_

   PIN u0_R2_26_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 6.706 0.163 6.734 ;
      END
   END u0_R2_26_

   PIN u0_R3_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.89 0.163 11.918 ;
      END
   END u0_R3_13_

   PIN u0_R3_16_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.338 0.0 52.366 0.163 ;
      END
   END u0_R3_16_

   PIN u0_R3_17_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.154 0.0 7.182 0.163 ;
      END
   END u0_R3_17_

   PIN u0_R3_19_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.73 0.163 15.758 ;
      END
   END u0_R3_19_

   PIN u0_R4_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.25 0.163 3.278 ;
      END
   END u0_R4_10_

   PIN u0_R4_17_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.922 0.163 23.95 ;
      END
   END u0_R4_17_

   PIN u0_R4_20_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.85 0.163 20.878 ;
      END
   END u0_R4_20_

   PIN u0_R5_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.97 94.557 17.998 94.72 ;
      END
   END u0_R5_13_

   PIN u0_R5_27_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.362 0.0 13.39 0.163 ;
      END
   END u0_R5_27_

   PIN u0_R5_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.386 94.557 6.414 94.72 ;
      END
   END u0_R5_4_

   PIN u0_R6_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.066 0.0 38.094 0.163 ;
      END
   END u0_R6_14_

   PIN u0_R6_17_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.794 0.163 15.822 ;
      END
   END u0_R6_17_

   PIN u0_R6_18_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.434 0.0 88.462 0.163 ;
      END
   END u0_R6_18_

   PIN u0_R6_23_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.274 0.0 100.302 0.163 ;
      END
   END u0_R6_23_

   PIN u0_R6_25_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.122 0.163 51.15 ;
      END
   END u0_R6_25_

   PIN u0_R6_26_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.426 0.0 117.454 0.163 ;
      END
   END u0_R6_26_

   PIN u0_R6_28_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.41 0.0 15.438 0.163 ;
      END
   END u0_R6_28_

   PIN u0_R6_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.146 0.0 20.174 0.163 ;
      END
   END u0_R6_3_

   PIN u0_R6_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.706 0.0 102.734 0.163 ;
      END
   END u0_R6_8_

   PIN u0_R7_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.498 0.0 64.526 0.163 ;
      END
   END u0_R7_10_

   PIN u0_R7_16_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.714 0.0 41.742 0.163 ;
      END
   END u0_R7_16_

   PIN u0_R7_20_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.09 0.0 63.118 0.163 ;
      END
   END u0_R7_20_

   PIN u0_R7_25_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.618 0.0 53.646 0.163 ;
      END
   END u0_R7_25_

   PIN u0_R7_28_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.578 0.0 38.606 0.163 ;
      END
   END u0_R7_28_

   PIN u0_R7_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.258 0.0 62.286 0.163 ;
      END
   END u0_R7_2_

   PIN u0_R7_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.818 0.0 40.846 0.163 ;
      END
   END u0_R7_6_

   PIN u0_R8_23_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.434 0.0 96.462 0.163 ;
      END
   END u0_R8_23_

   PIN u0_key_r_23_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.786 0.0 36.814 0.163 ;
      END
   END u0_key_r_23_

   PIN u0_key_r_44_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.938 0.0 5.966 0.163 ;
      END
   END u0_key_r_44_

   PIN u0_uk_K_r_251
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.002 0.0 6.03 0.163 ;
      END
   END u0_uk_K_r_251

   PIN u0_uk_K_r_263
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.05 0.163 8.078 ;
      END
   END u0_uk_K_r_263

   PIN u0_uk_K_r_273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.282 0.0 7.31 0.163 ;
      END
   END u0_uk_K_r_273

   PIN u0_uk_K_r_332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.738 0.163 10.766 ;
      END
   END u0_uk_K_r_332

   PIN u0_uk_K_r_335
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.394 0.0 1.422 0.163 ;
      END
   END u0_uk_K_r_335

   PIN u0_uk_K_r_343
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.522 0.0 1.55 0.163 ;
      END
   END u0_uk_K_r_343

   PIN u0_uk_K_r_344
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.626 0.0 0.654 0.163 ;
      END
   END u0_uk_K_r_344

   PIN u0_uk_K_r_356
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.418 0.0 2.446 0.163 ;
      END
   END u0_uk_K_r_356

   PIN u0_uk_K_r_357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.114 0.163 24.142 ;
      END
   END u0_uk_K_r_357

   PIN u0_uk_K_r_359
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.954 0.163 19.982 ;
      END
   END u0_uk_K_r_359

   PIN u0_uk_K_r_365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.562 0.0 0.59 0.163 ;
      END
   END u0_uk_K_r_365

   PIN u0_uk_K_r_378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.354 0.0 2.382 0.163 ;
      END
   END u0_uk_K_r_378

   PIN u0_uk_K_r_381
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.49 0.0 5.518 0.163 ;
      END
   END u0_uk_K_r_381

   PIN u0_uk_K_r_401
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.026 0.163 7.054 ;
      END
   END u0_uk_K_r_401

   PIN u0_uk_K_r_413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.61 0.163 10.638 ;
      END
   END u0_uk_K_r_413

   PIN u0_uk_K_r_437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.33 0.0 1.358 0.163 ;
      END
   END u0_uk_K_r_437

   PIN u0_uk_K_r_449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.338 0.0 4.366 0.163 ;
      END
   END u0_uk_K_r_449

   PIN u0_uk_K_r_530
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.738 0.0 10.766 0.163 ;
      END
   END u0_uk_K_r_530

   PIN u1_L10_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.914 0.0 12.942 0.163 ;
      END
   END u1_L10_13_

   PIN u1_L11_22_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.826 0.163 11.854 ;
      END
   END u1_L11_22_

   PIN u1_L11_reg_7__Q
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.218 0.163 15.246 ;
      END
   END u1_L11_reg_7__Q

   PIN u1_L7_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.698 0.163 11.726 ;
      END
   END u1_L7_7_

   PIN u1_R10_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.17 0.163 13.198 ;
      END
   END u1_R10_12_

   PIN u1_R8_19_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.106 0.163 13.134 ;
      END
   END u1_R8_19_

   PIN u1_R8_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.778 94.557 17.806 94.72 ;
      END
   END u1_R8_7_

   PIN u2_R6_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.866 0.0 98.894 0.163 ;
      END
   END u2_R6_7_

   PIN u2_R7_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.29 0.0 74.318 0.163 ;
      END
   END u2_R7_15_

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 175.744 94.72 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 175.744 94.72 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 175.744 94.72 ;
      LAYER V1 ;
         RECT 0.0 0.0 175.744 94.72 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 175.744 94.72 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 175.744 94.72 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 175.744 94.72 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 175.744 94.72 ;
      LAYER M1 ;
         RECT 0.0 0.0 175.744 94.72 ;
   END
END h3_mgc_des_perf_a

MACRO h2_mgc_des_perf_a
   CLASS BLOCK ;
   FOREIGN h2 ;
   ORIGIN 0 0 ;
   SIZE 167.36 BY 61.44 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1114_n_21429
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.57 61.277 51.598 61.44 ;
      END
   END FE_OFN1114_n_21429

   PIN FE_OFN1152_n_14527
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.234 61.277 93.262 61.44 ;
      END
   END FE_OFN1152_n_14527

   PIN FE_OFN1308_n_14014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.442 61.277 67.47 61.44 ;
      END
   END FE_OFN1308_n_14014

   PIN FE_OFN13_n_106596
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.37 0.0 64.398 0.163 ;
      END
   END FE_OFN13_n_106596

   PIN FE_OFN1911_n_80620
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.138 61.277 33.166 61.44 ;
      END
   END FE_OFN1911_n_80620

   PIN FE_OFN194_n_84781
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.01 61.277 33.038 61.44 ;
      END
   END FE_OFN194_n_84781

   PIN FE_OFN200_n_15151
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.466 61.277 52.494 61.44 ;
      END
   END FE_OFN200_n_15151

   PIN FE_OFN2035_n_14525
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.234 61.277 53.262 61.44 ;
      END
   END FE_OFN2035_n_14525

   PIN FE_OFN2064_g190297_u0_o
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 157.426 61.277 157.454 61.44 ;
      END
   END FE_OFN2064_g190297_u0_o

   PIN FE_OFN2073_n_107830
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.402 0.0 156.43 0.163 ;
      END
   END FE_OFN2073_n_107830

   PIN FE_OFN2234_n_75724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.434 61.277 32.462 61.44 ;
      END
   END FE_OFN2234_n_75724

   PIN FE_OFN2250_n_82961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.058 61.277 83.086 61.44 ;
      END
   END FE_OFN2250_n_82961

   PIN FE_OFN22_n_104304
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.274 61.277 92.302 61.44 ;
      END
   END FE_OFN22_n_104304

   PIN FE_OFN245_n_79557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.922 61.277 63.95 61.44 ;
      END
   END FE_OFN245_n_79557

   PIN FE_OFN2549_n_118022
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.826 61.277 147.854 61.44 ;
      END
   END FE_OFN2549_n_118022

   PIN FE_OFN2763_n_107068
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.458 61.277 153.486 61.44 ;
      END
   END FE_OFN2763_n_107068

   PIN FE_OFN3492_n_83012
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.378 61.277 75.406 61.44 ;
      END
   END FE_OFN3492_n_83012

   PIN FE_OFN3552_n_81000
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.314 61.277 59.342 61.44 ;
      END
   END FE_OFN3552_n_81000

   PIN FE_OFN3554_n_108480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 59.186 167.36 59.214 ;
      END
   END FE_OFN3554_n_108480

   PIN FE_OFN4785_n_77924
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.754 61.277 8.782 61.44 ;
      END
   END FE_OFN4785_n_77924

   PIN FE_OFN818_n_103115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.762 61.277 75.79 61.44 ;
      END
   END FE_OFN818_n_103115

   PIN FE_OFN867_n_14026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.17 61.277 37.198 61.44 ;
      END
   END FE_OFN867_n_14026

   PIN desOut_16_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.458 0.0 129.486 0.163 ;
      END
   END desOut_16_

   PIN desOut_17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.818 0.0 144.846 0.163 ;
      END
   END desOut_17_

   PIN desOut_38_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.138 0.0 41.166 0.163 ;
      END
   END desOut_38_

   PIN g190280_u0_o
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.178 0.0 160.206 0.163 ;
      END
   END g190280_u0_o

   PIN g190611_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 147.89 61.277 147.918 61.44 ;
      END
   END g190611_p

   PIN g190906_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 15.282 167.36 15.31 ;
      END
   END g190906_p

   PIN g190953_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 49.522 167.36 49.55 ;
      END
   END g190953_p

   PIN g191131_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 49.778 167.36 49.806 ;
      END
   END g191131_p

   PIN g191163_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 49.586 167.36 49.614 ;
      END
   END g191163_p

   PIN g191647_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.714 61.277 121.742 61.44 ;
      END
   END g191647_da

   PIN g191647_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.178 61.277 120.206 61.44 ;
      END
   END g191647_db

   PIN g191648_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.146 0.0 52.174 0.163 ;
      END
   END g191648_da

   PIN g191648_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.154 0.0 55.182 0.163 ;
      END
   END g191648_db

   PIN g192426_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.61 61.277 114.638 61.44 ;
      END
   END g192426_p

   PIN g192601_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.018 61.277 60.046 61.44 ;
      END
   END g192601_p

   PIN g192862_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.162 0.163 26.19 ;
      END
   END g192862_p

   PIN g192893_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.706 0.163 22.734 ;
      END
   END g192893_p

   PIN g193052_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.858 0.0 71.886 0.163 ;
      END
   END g193052_p

   PIN g195141_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.114 61.277 48.142 61.44 ;
      END
   END g195141_da

   PIN g195175_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.546 61.277 90.574 61.44 ;
      END
   END g195175_p

   PIN g218222_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.17 61.277 93.198 61.44 ;
      END
   END g218222_sb

   PIN g218659_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.346 61.277 55.374 61.44 ;
      END
   END g218659_da

   PIN g218659_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.97 61.277 57.998 61.44 ;
      END
   END g218659_db

   PIN g219318_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.546 61.277 98.574 61.44 ;
      END
   END g219318_p

   PIN g219362_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.466 61.277 28.494 61.44 ;
      END
   END g219362_p

   PIN g219365_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.562 61.277 96.59 61.44 ;
      END
   END g219365_p

   PIN g220459_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.298 61.277 29.326 61.44 ;
      END
   END g220459_da

   PIN g220459_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.106 61.277 29.134 61.44 ;
      END
   END g220459_db

   PIN g223661_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.858 61.277 39.886 61.44 ;
      END
   END g223661_p

   PIN g223834_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.93 61.277 34.958 61.44 ;
      END
   END g223834_sb

   PIN g288188_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.626 61.277 72.654 61.44 ;
      END
   END g288188_p

   PIN g288202_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.554 61.277 69.582 61.44 ;
      END
   END g288202_p

   PIN g288612_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.458 61.277 25.486 61.44 ;
      END
   END g288612_p

   PIN key_c_r_31__2158
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.386 61.277 70.414 61.44 ;
      END
   END key_c_r_31__2158

   PIN key_c_r_33__8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.186 61.277 83.214 61.44 ;
      END
   END key_c_r_33__8_

   PIN n_100862
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.13 61.277 110.158 61.44 ;
      END
   END n_100862

   PIN n_100928
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.722 0.0 116.75 0.163 ;
      END
   END n_100928

   PIN n_101021
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 136.882 61.277 136.91 61.44 ;
      END
   END n_101021

   PIN n_102321
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 133.362 61.277 133.39 61.44 ;
      END
   END n_102321

   PIN n_102578
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 130.994 61.277 131.022 61.44 ;
      END
   END n_102578

   PIN n_103024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 156.402 61.277 156.43 61.44 ;
      END
   END n_103024

   PIN n_103133
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.058 61.277 83.086 61.44 ;
      END
   END n_103133

   PIN n_103323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.65 61.358 89.678 61.44 ;
      END
   END n_103323

   PIN n_103421
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.378 61.277 83.406 61.44 ;
      END
   END n_103421

   PIN n_103511
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.362 61.277 93.39 61.44 ;
      END
   END n_103511

   PIN n_103611
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.674 61.277 90.702 61.44 ;
      END
   END n_103611

   PIN n_103663
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.498 61.277 88.526 61.44 ;
      END
   END n_103663

   PIN n_103665
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.082 61.277 92.11 61.44 ;
      END
   END n_103665

   PIN n_103666
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.114 61.277 88.142 61.44 ;
      END
   END n_103666

   PIN n_103777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.514 61.277 78.542 61.44 ;
      END
   END n_103777

   PIN n_103800
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.738 61.277 90.766 61.44 ;
      END
   END n_103800

   PIN n_103935
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.674 61.277 90.702 61.44 ;
      END
   END n_103935

   PIN n_104032
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.81 61.277 85.838 61.44 ;
      END
   END n_104032

   PIN n_104077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.09 61.277 79.118 61.44 ;
      END
   END n_104077

   PIN n_104097
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.69 61.277 88.718 61.44 ;
      END
   END n_104097

   PIN n_104144
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.962 61.277 86.99 61.44 ;
      END
   END n_104144

   PIN n_104146
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.13 61.277 78.158 61.44 ;
      END
   END n_104146

   PIN n_104171
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.122 61.277 83.15 61.44 ;
      END
   END n_104171

   PIN n_104175
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.25 61.277 83.278 61.44 ;
      END
   END n_104175

   PIN n_104263
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.57 61.277 83.598 61.44 ;
      END
   END n_104263

   PIN n_104285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.074 61.277 81.102 61.44 ;
      END
   END n_104285

   PIN n_104385
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.442 61.277 83.47 61.44 ;
      END
   END n_104385

   PIN n_104389
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.178 61.277 88.206 61.44 ;
      END
   END n_104389

   PIN n_104484
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.506 61.277 99.534 61.44 ;
      END
   END n_104484

   PIN n_104500
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.194 61.277 78.222 61.44 ;
      END
   END n_104500

   PIN n_104533
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 84.978 61.277 85.006 61.44 ;
      END
   END n_104533

   PIN n_104591
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.13 61.277 78.158 61.44 ;
      END
   END n_104591

   PIN n_104636
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.426 61.277 85.454 61.44 ;
      END
   END n_104636

   PIN n_104655
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.442 61.277 75.47 61.44 ;
      END
   END n_104655

   PIN n_104669
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.29 61.277 74.318 61.44 ;
      END
   END n_104669

   PIN n_105032
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.426 0.0 77.454 0.163 ;
      END
   END n_105032

   PIN n_105114
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.986 0.0 72.014 0.082 ;
      END
   END n_105114

   PIN n_105153
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.786 61.277 52.814 61.44 ;
      END
   END n_105153

   PIN n_105173
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.21 0.0 68.238 0.163 ;
      END
   END n_105173

   PIN n_105210
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.97 0.163 25.998 ;
      END
   END n_105210

   PIN n_105221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.546 0.163 26.574 ;
      END
   END n_105221

   PIN n_105285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.002 0.163 22.03 ;
      END
   END n_105285

   PIN n_105324
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.746 61.277 125.774 61.44 ;
      END
   END n_105324

   PIN n_105338
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.226 0.163 26.254 ;
      END
   END n_105338

   PIN n_105358
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.506 0.163 35.534 ;
      END
   END n_105358

   PIN n_105422
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.666 0.0 71.694 0.163 ;
      END
   END n_105422

   PIN n_105473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.674 61.277 114.702 61.44 ;
      END
   END n_105473

   PIN n_105532
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.386 0.163 30.414 ;
      END
   END n_105532

   PIN n_105558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.41 0.0 79.438 0.163 ;
      END
   END n_105558

   PIN n_105559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.05 0.0 64.078 0.163 ;
      END
   END n_105559

   PIN n_105594
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.602 0.0 79.63 0.163 ;
      END
   END n_105594

   PIN n_105646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.986 0.0 64.014 0.163 ;
      END
   END n_105646

   PIN n_105647
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.786 0.0 68.814 0.163 ;
      END
   END n_105647

   PIN n_105690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.658 0.0 52.686 0.163 ;
      END
   END n_105690

   PIN n_105698
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.386 61.277 118.414 61.44 ;
      END
   END n_105698

   PIN n_105744
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.89 0.0 67.918 0.163 ;
      END
   END n_105744

   PIN n_105750
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.146 0.0 60.174 0.163 ;
      END
   END n_105750

   PIN n_105751
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.538 0.0 79.566 0.163 ;
      END
   END n_105751

   PIN n_105789
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.754 0.163 16.782 ;
      END
   END n_105789

   PIN n_105899
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 19.122 0.163 19.15 ;
      END
   END n_105899

   PIN n_105911
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.21 0.0 60.238 0.163 ;
      END
   END n_105911

   PIN n_105913
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.498 0.0 56.526 0.163 ;
      END
   END n_105913

   PIN n_105936
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.97 0.0 57.998 0.163 ;
      END
   END n_105936

   PIN n_105940
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.49 0.0 77.518 0.082 ;
      END
   END n_105940

   PIN n_105951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.506 0.163 19.534 ;
      END
   END n_105951

   PIN n_105999
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.322 61.277 118.35 61.44 ;
      END
   END n_105999

   PIN n_106024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.202 61.277 113.23 61.44 ;
      END
   END n_106024

   PIN n_106031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.754 0.0 48.782 0.163 ;
      END
   END n_106031

   PIN n_106032
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.178 0.0 64.206 0.163 ;
      END
   END n_106032

   PIN n_106044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.082 61.277 124.11 61.44 ;
      END
   END n_106044

   PIN n_106048
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.738 0.0 98.766 0.163 ;
      END
   END n_106048

   PIN n_106077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.186 0.163 19.214 ;
      END
   END n_106077

   PIN n_106100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.77 0.163 22.798 ;
      END
   END n_106100

   PIN n_106152
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.698 0.163 19.726 ;
      END
   END n_106152

   PIN n_106178
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.81 0.163 21.838 ;
      END
   END n_106178

   PIN n_106206
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.85 61.277 116.878 61.44 ;
      END
   END n_106206

   PIN n_106225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.018 0.0 60.046 0.163 ;
      END
   END n_106225

   PIN n_106257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.57 0.163 19.598 ;
      END
   END n_106257

   PIN n_106305
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.242 61.277 120.27 61.44 ;
      END
   END n_106305

   PIN n_106309
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.37 61.277 120.398 61.44 ;
      END
   END n_106309

   PIN n_106315
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.362 0.0 61.39 0.163 ;
      END
   END n_106315

   PIN n_106345
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.65 61.277 121.678 61.44 ;
      END
   END n_106345

   PIN n_106356
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.282 0.0 63.31 0.163 ;
      END
   END n_106356

   PIN n_106374
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.842 0.163 25.87 ;
      END
   END n_106374

   PIN n_106382
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 165.362 61.277 165.39 61.44 ;
      END
   END n_106382

   PIN n_106401
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.122 61.277 123.15 61.44 ;
      END
   END n_106401

   PIN n_106404
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.514 0.163 30.542 ;
      END
   END n_106404

   PIN n_106446
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.722 0.0 52.75 0.163 ;
      END
   END n_106446

   PIN n_106447
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.818 0.0 48.846 0.163 ;
      END
   END n_106447

   PIN n_106458
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.026 0.163 15.054 ;
      END
   END n_106458

   PIN n_106496
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.586 61.277 121.614 61.44 ;
      END
   END n_106496

   PIN n_106527
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.874 0.163 21.902 ;
      END
   END n_106527

   PIN n_106534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.562 0.163 16.59 ;
      END
   END n_106534

   PIN n_106558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.938 0.0 37.966 0.163 ;
      END
   END n_106558

   PIN n_106576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.634 0.163 19.662 ;
      END
   END n_106576

   PIN n_106582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.362 0.163 21.39 ;
      END
   END n_106582

   PIN n_106653
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.522 61.277 121.55 61.44 ;
      END
   END n_106653

   PIN n_106665
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.466 0.0 52.494 0.163 ;
      END
   END n_106665

   PIN n_106667
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.818 0.163 16.846 ;
      END
   END n_106667

   PIN n_106671
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.986 61.277 64.014 61.44 ;
      END
   END n_106671

   PIN n_106682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.674 61.277 122.702 61.44 ;
      END
   END n_106682

   PIN n_106715
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.602 0.0 39.63 0.163 ;
      END
   END n_106715

   PIN n_106742
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.682 61.277 125.71 61.44 ;
      END
   END n_106742

   PIN n_106753
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.474 61.277 71.502 61.44 ;
      END
   END n_106753

   PIN n_106769
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.418 61.277 42.446 61.44 ;
      END
   END n_106769

   PIN n_106772
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.082 61.277 60.11 61.44 ;
      END
   END n_106772

   PIN n_106806
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.69 61.277 144.718 61.44 ;
      END
   END n_106806

   PIN n_106814
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.498 0.0 48.526 0.163 ;
      END
   END n_106814

   PIN n_106816
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.362 0.0 45.39 0.163 ;
      END
   END n_106816

   PIN n_106875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.274 61.277 52.302 61.44 ;
      END
   END n_106875

   PIN n_107039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.306 61.277 160.334 61.44 ;
      END
   END n_107039

   PIN n_107087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.57 0.0 163.598 0.163 ;
      END
   END n_107087

   PIN n_107115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 53.682 167.36 53.71 ;
      END
   END n_107115

   PIN n_107137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.146 61.277 164.174 61.44 ;
      END
   END n_107137

   PIN n_107138
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.786 61.277 148.814 61.44 ;
      END
   END n_107138

   PIN n_107156
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.018 61.277 164.046 61.44 ;
      END
   END n_107156

   PIN n_107223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.178 61.277 152.206 61.44 ;
      END
   END n_107223

   PIN n_107261
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 148.466 61.277 148.494 61.44 ;
      END
   END n_107261

   PIN n_107361
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.082 61.277 164.11 61.44 ;
      END
   END n_107361

   PIN n_107390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.69 61.277 152.718 61.44 ;
      END
   END n_107390

   PIN n_107391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.242 61.277 152.27 61.44 ;
      END
   END n_107391

   PIN n_107409
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.73 0.0 159.758 0.163 ;
      END
   END n_107409

   PIN n_107414
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 148.594 61.277 148.622 61.44 ;
      END
   END n_107414

   PIN n_107424
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 163.058 0.0 163.086 0.163 ;
      END
   END n_107424

   PIN n_107426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.626 0.0 144.654 0.163 ;
      END
   END n_107426

   PIN n_107429
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 11.762 167.36 11.79 ;
      END
   END n_107429

   PIN n_107430
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.114 0.0 160.142 0.163 ;
      END
   END n_107430

   PIN n_107482
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 148.658 61.277 148.686 61.44 ;
      END
   END n_107482

   PIN n_107485
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 45.938 167.36 45.966 ;
      END
   END n_107485

   PIN n_107498
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.018 0.0 164.046 0.163 ;
      END
   END n_107498

   PIN n_107515
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 148.722 61.277 148.75 61.44 ;
      END
   END n_107515

   PIN n_107520
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.146 61.277 156.174 61.44 ;
      END
   END n_107520

   PIN n_107556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 25.97 167.36 25.998 ;
      END
   END n_107556

   PIN n_107586
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 3.762 167.36 3.79 ;
      END
   END n_107586

   PIN n_107658
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.242 0.0 160.27 0.163 ;
      END
   END n_107658

   PIN n_107704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 25.842 167.36 25.87 ;
      END
   END n_107704

   PIN n_107733
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.178 61.277 160.206 61.44 ;
      END
   END n_107733

   PIN n_107740
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.554 0.0 125.582 0.163 ;
      END
   END n_107740

   PIN n_107831
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.25 0.0 163.278 0.163 ;
      END
   END n_107831

   PIN n_107875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.594 61.277 148.622 61.44 ;
      END
   END n_107875

   PIN n_107879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 158.898 0.0 158.926 0.163 ;
      END
   END n_107879

   PIN n_107901
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.498 0.0 152.526 0.163 ;
      END
   END n_107901

   PIN n_107909
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.434 61.277 152.462 61.44 ;
      END
   END n_107909

   PIN n_107910
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.13 0.0 150.158 0.163 ;
      END
   END n_107910

   PIN n_107929
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 160.178 61.277 160.206 61.44 ;
      END
   END n_107929

   PIN n_107930
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.106 61.277 149.134 61.44 ;
      END
   END n_107930

   PIN n_107938
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 154.738 61.277 154.766 61.44 ;
      END
   END n_107938

   PIN n_107997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.274 61.277 156.302 61.44 ;
      END
   END n_107997

   PIN n_107998
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.562 0.0 144.59 0.163 ;
      END
   END n_107998

   PIN n_108000
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 38.322 167.36 38.35 ;
      END
   END n_108000

   PIN n_108052
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.21 61.277 164.238 61.44 ;
      END
   END n_108052

   PIN n_108056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 156.082 61.358 156.11 61.44 ;
      END
   END n_108056

   PIN n_108058
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 148.53 61.277 148.558 61.44 ;
      END
   END n_108058

   PIN n_108059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 148.402 61.277 148.43 61.44 ;
      END
   END n_108059

   PIN n_108064
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.138 0.0 161.166 0.163 ;
      END
   END n_108064

   PIN n_108065
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 26.674 167.36 26.702 ;
      END
   END n_108065

   PIN n_108083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.186 61.277 147.214 61.44 ;
      END
   END n_108083

   PIN n_108088
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.338 0.0 156.366 0.163 ;
      END
   END n_108088

   PIN n_108129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 16.242 167.36 16.27 ;
      END
   END n_108129

   PIN n_108132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.818 0.0 160.846 0.163 ;
      END
   END n_108132

   PIN n_108133
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 149.554 0.0 149.582 0.163 ;
      END
   END n_108133

   PIN n_108161
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.114 61.277 152.142 61.44 ;
      END
   END n_108161

   PIN n_108172
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.626 61.277 152.654 61.44 ;
      END
   END n_108172

   PIN n_108179
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.41 61.277 143.438 61.44 ;
      END
   END n_108179

   PIN n_108192
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.962 61.277 142.99 61.44 ;
      END
   END n_108192

   PIN n_108216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 23.026 167.36 23.054 ;
      END
   END n_108216

   PIN n_108224
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.242 61.277 160.27 61.44 ;
      END
   END n_108224

   PIN n_108227
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 26.802 167.36 26.83 ;
      END
   END n_108227

   PIN n_108234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.562 61.277 152.59 61.44 ;
      END
   END n_108234

   PIN n_108235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.498 61.277 152.526 61.44 ;
      END
   END n_108235

   PIN n_108244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 39.986 167.36 40.014 ;
      END
   END n_108244

   PIN n_108274
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.274 61.277 164.302 61.44 ;
      END
   END n_108274

   PIN n_108297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 59.122 167.36 59.15 ;
      END
   END n_108297

   PIN n_108300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.562 61.277 152.59 61.44 ;
      END
   END n_108300

   PIN n_108311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.306 61.277 152.334 61.44 ;
      END
   END n_108311

   PIN n_108318
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.754 61.277 152.782 61.44 ;
      END
   END n_108318

   PIN n_108320
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.754 61.277 152.782 61.44 ;
      END
   END n_108320

   PIN n_108329
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.626 61.277 152.654 61.44 ;
      END
   END n_108329

   PIN n_108337
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 59.25 167.36 59.278 ;
      END
   END n_108337

   PIN n_108392
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 49.65 167.36 49.678 ;
      END
   END n_108392

   PIN n_108450
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.818 61.277 152.846 61.44 ;
      END
   END n_108450

   PIN n_108486
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.986 61.277 152.014 61.44 ;
      END
   END n_108486

   PIN n_112858
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.73 61.277 79.758 61.44 ;
      END
   END n_112858

   PIN n_112987
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.018 0.0 148.046 0.163 ;
      END
   END n_112987

   PIN n_117115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.842 61.277 81.87 61.44 ;
      END
   END n_117115

   PIN n_118365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.21 61.277 92.238 61.44 ;
      END
   END n_118365

   PIN n_118376
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.754 61.277 88.782 61.44 ;
      END
   END n_118376

   PIN n_118637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.65 61.277 121.678 61.44 ;
      END
   END n_118637

   PIN n_126056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.954 61.277 107.982 61.44 ;
      END
   END n_126056

   PIN n_126215
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.762 0.163 11.79 ;
      END
   END n_126215

   PIN n_13159
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.786 61.277 44.814 61.44 ;
      END
   END n_13159

   PIN n_13183
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.618 61.277 37.646 61.44 ;
      END
   END n_13183

   PIN n_13379
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.298 61.277 29.326 61.44 ;
      END
   END n_13379

   PIN n_13383
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.45 61.277 46.478 61.44 ;
      END
   END n_13383

   PIN n_13413
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.666 61.277 71.694 61.44 ;
      END
   END n_13413

   PIN n_13426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.01 61.277 33.038 61.44 ;
      END
   END n_13426

   PIN n_13478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.594 61.277 28.622 61.44 ;
      END
   END n_13478

   PIN n_13607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.826 61.277 35.854 61.44 ;
      END
   END n_13607

   PIN n_13698
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.426 61.277 37.454 61.44 ;
      END
   END n_13698

   PIN n_137144
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.602 0.163 7.63 ;
      END
   END n_137144

   PIN n_137150
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.826 0.163 11.854 ;
      END
   END n_137150

   PIN n_13862
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.282 61.277 47.31 61.44 ;
      END
   END n_13862

   PIN n_13873
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.962 61.277 70.99 61.44 ;
      END
   END n_13873

   PIN n_13932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.546 61.277 66.574 61.44 ;
      END
   END n_13932

   PIN n_14044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.698 61.277 67.726 61.44 ;
      END
   END n_14044

   PIN n_14147
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.282 61.277 63.31 61.44 ;
      END
   END n_14147

   PIN n_14374
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.226 61.277 50.254 61.44 ;
      END
   END n_14374

   PIN n_14380
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.178 61.277 48.206 61.44 ;
      END
   END n_14380

   PIN n_183945
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.394 61.277 33.422 61.44 ;
      END
   END n_183945

   PIN n_183950
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 21.362 167.36 21.39 ;
      END
   END n_183950

   PIN n_75398
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.41 61.277 39.438 61.44 ;
      END
   END n_75398

   PIN n_75503
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.098 61.277 34.126 61.44 ;
      END
   END n_75503

   PIN n_75797
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.522 61.277 25.55 61.44 ;
      END
   END n_75797

   PIN n_75845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.778 61.277 25.806 61.44 ;
      END
   END n_75845

   PIN n_75864
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.61 61.277 90.638 61.44 ;
      END
   END n_75864

   PIN n_75994
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.002 61.277 38.03 61.44 ;
      END
   END n_75994

   PIN n_76007
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.562 61.277 160.59 61.44 ;
      END
   END n_76007

   PIN n_76135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.426 61.277 21.454 61.44 ;
      END
   END n_76135

   PIN n_76204
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.554 61.277 37.582 61.44 ;
      END
   END n_76204

   PIN n_76218
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.05 61.277 64.078 61.44 ;
      END
   END n_76218

   PIN n_76344
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.202 61.277 129.23 61.44 ;
      END
   END n_76344

   PIN n_76528
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.682 61.277 21.71 61.44 ;
      END
   END n_76528

   PIN n_76756
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.642 61.277 14.67 61.44 ;
      END
   END n_76756

   PIN n_76912
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.426 61.277 13.454 61.44 ;
      END
   END n_76912

   PIN n_76917
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.074 61.277 25.102 61.44 ;
      END
   END n_76917

   PIN n_76933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.146 61.277 20.174 61.44 ;
      END
   END n_76933

   PIN n_76936
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.194 61.277 6.222 61.44 ;
      END
   END n_76936

   PIN n_76947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.746 61.277 21.774 61.44 ;
      END
   END n_76947

   PIN n_76948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.122 61.277 27.15 61.44 ;
      END
   END n_76948

   PIN n_76988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.098 61.277 18.126 61.44 ;
      END
   END n_76988

   PIN n_77102
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.514 61.277 14.542 61.44 ;
      END
   END n_77102

   PIN n_77104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.882 61.277 0.91 61.44 ;
      END
   END n_77104

   PIN n_77105
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.418 61.277 10.446 61.44 ;
      END
   END n_77105

   PIN n_77161
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.226 61.277 10.254 61.44 ;
      END
   END n_77161

   PIN n_77283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.946 61.277 0.974 61.44 ;
      END
   END n_77283

   PIN n_77379
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.05 61.277 16.078 61.44 ;
      END
   END n_77379

   PIN n_77468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.226 61.277 10.254 61.44 ;
      END
   END n_77468

   PIN n_77547
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.29 61.277 2.318 61.44 ;
      END
   END n_77547

   PIN n_77747
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.13 61.277 14.158 61.44 ;
      END
   END n_77747

   PIN n_77781
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.482 61.277 10.51 61.44 ;
      END
   END n_77781

   PIN n_77819
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.29 61.277 10.318 61.44 ;
      END
   END n_77819

   PIN n_78099
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.602 61.277 7.63 61.44 ;
      END
   END n_78099

   PIN n_78517
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.17 61.277 5.198 61.44 ;
      END
   END n_78517

   PIN n_78714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.25 61.277 27.278 61.44 ;
      END
   END n_78714

   PIN n_78796
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.578 61.277 22.606 61.44 ;
      END
   END n_78796

   PIN n_78872
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.898 61.277 22.926 61.44 ;
      END
   END n_78872

   PIN n_78903
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.442 61.277 59.47 61.44 ;
      END
   END n_78903

   PIN n_78996
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.538 61.277 71.566 61.44 ;
      END
   END n_78996

   PIN n_79015
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.786 61.277 132.814 61.44 ;
      END
   END n_79015

   PIN n_79054
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.986 61.277 136.014 61.44 ;
      END
   END n_79054

   PIN n_79058
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.106 61.277 133.134 61.44 ;
      END
   END n_79058

   PIN n_79069
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.954 61.277 75.982 61.44 ;
      END
   END n_79069

   PIN n_79114
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.218 61.277 31.246 61.44 ;
      END
   END n_79114

   PIN n_79207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.826 61.358 107.854 61.44 ;
      END
   END n_79207

   PIN n_79217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.53 61.277 140.558 61.44 ;
      END
   END n_79217

   PIN n_79224
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 140.978 61.277 141.006 61.44 ;
      END
   END n_79224

   PIN n_79290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.554 61.277 37.582 61.44 ;
      END
   END n_79290

   PIN n_79306
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.81 61.358 37.838 61.44 ;
      END
   END n_79306

   PIN n_79355
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.162 61.277 138.19 61.44 ;
      END
   END n_79355

   PIN n_79357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 137.01 61.277 137.038 61.44 ;
      END
   END n_79357

   PIN n_79378
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 140.402 61.277 140.43 61.44 ;
      END
   END n_79378

   PIN n_79379
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 141.618 61.277 141.646 61.44 ;
      END
   END n_79379

   PIN n_79388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.162 61.277 58.19 61.44 ;
      END
   END n_79388

   PIN n_79399
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.218 61.277 135.246 61.44 ;
      END
   END n_79399

   PIN n_79410
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.202 61.277 33.23 61.44 ;
      END
   END n_79410

   PIN n_79432
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.186 61.277 107.214 61.44 ;
      END
   END n_79432

   PIN n_79456
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.586 61.277 33.614 61.44 ;
      END
   END n_79456

   PIN n_79462
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.658 61.277 140.686 61.44 ;
      END
   END n_79462

   PIN n_79483
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.146 61.277 132.174 61.44 ;
      END
   END n_79483

   PIN n_79497
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.538 61.277 79.566 61.44 ;
      END
   END n_79497

   PIN n_79507
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.626 61.277 48.654 61.44 ;
      END
   END n_79507

   PIN n_79513
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.202 61.358 41.23 61.44 ;
      END
   END n_79513

   PIN n_79516
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 57.33 61.277 57.358 61.44 ;
      END
   END n_79516

   PIN n_79537
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.85 61.277 44.878 61.44 ;
      END
   END n_79537

   PIN n_79569
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.058 61.277 59.086 61.44 ;
      END
   END n_79569

   PIN n_79577
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.41 61.358 47.438 61.44 ;
      END
   END n_79577

   PIN n_79626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.178 61.277 64.206 61.44 ;
      END
   END n_79626

   PIN n_79648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.498 61.358 88.526 61.44 ;
      END
   END n_79648

   PIN n_79650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 129.266 61.277 129.294 61.44 ;
      END
   END n_79650

   PIN n_79680
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.082 61.277 76.11 61.44 ;
      END
   END n_79680

   PIN n_79682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.818 61.277 40.846 61.44 ;
      END
   END n_79682

   PIN n_79688
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.69 61.277 56.718 61.44 ;
      END
   END n_79688

   PIN n_79690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.866 61.277 34.894 61.44 ;
      END
   END n_79690

   PIN n_79712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.042 61.277 133.07 61.44 ;
      END
   END n_79712

   PIN n_79715
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.266 61.277 33.294 61.44 ;
      END
   END n_79715

   PIN n_79718
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.578 0.0 110.606 0.163 ;
      END
   END n_79718

   PIN n_79779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.954 61.277 139.982 61.44 ;
      END
   END n_79779

   PIN n_79782
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 136.818 61.277 136.846 61.44 ;
      END
   END n_79782

   PIN n_79783
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.978 61.277 133.006 61.44 ;
      END
   END n_79783

   PIN n_79785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 135.346 61.277 135.374 61.44 ;
      END
   END n_79785

   PIN n_79863
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.154 61.277 79.182 61.44 ;
      END
   END n_79863

   PIN n_79879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.426 61.277 29.454 61.44 ;
      END
   END n_79879

   PIN n_79888
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.85 61.277 52.878 61.44 ;
      END
   END n_79888

   PIN n_79920
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 133.298 61.277 133.326 61.44 ;
      END
   END n_79920

   PIN n_79923
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.49 61.277 133.518 61.44 ;
      END
   END n_79923

   PIN n_79934
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 137.074 61.277 137.102 61.44 ;
      END
   END n_79934

   PIN n_79946
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.146 61.277 60.174 61.44 ;
      END
   END n_79946

   PIN n_79982
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.81 0.0 93.838 0.163 ;
      END
   END n_79982

   PIN n_79989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.466 61.277 108.494 61.44 ;
      END
   END n_79989

   PIN n_80001
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.554 61.277 45.582 61.44 ;
      END
   END n_80001

   PIN n_80015
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.314 61.277 91.342 61.44 ;
      END
   END n_80015

   PIN n_80058
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.762 61.277 139.79 61.44 ;
      END
   END n_80058

   PIN n_80061
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.77 61.277 142.798 61.44 ;
      END
   END n_80061

   PIN n_80062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.426 61.277 133.454 61.44 ;
      END
   END n_80062

   PIN n_80214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.882 61.277 136.91 61.44 ;
      END
   END n_80214

   PIN n_80220
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.61 61.277 90.638 61.44 ;
      END
   END n_80220

   PIN n_80221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.218 61.277 79.246 61.44 ;
      END
   END n_80221

   PIN n_80223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.834 0.0 94.862 0.163 ;
      END
   END n_80223

   PIN n_80226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.754 61.277 136.782 61.44 ;
      END
   END n_80226

   PIN n_80246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.946 61.277 136.974 61.44 ;
      END
   END n_80246

   PIN n_80251
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.914 61.277 44.942 61.44 ;
      END
   END n_80251

   PIN n_80267
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.522 61.277 33.55 61.44 ;
      END
   END n_80267

   PIN n_80270
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.546 61.277 130.574 61.44 ;
      END
   END n_80270

   PIN n_80310
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.33 61.277 33.358 61.44 ;
      END
   END n_80310

   PIN n_80338
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 137.138 61.277 137.166 61.44 ;
      END
   END n_80338

   PIN n_80339
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.722 61.277 140.75 61.44 ;
      END
   END n_80339

   PIN n_80391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.882 61.277 40.91 61.44 ;
      END
   END n_80391

   PIN n_80400
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.522 61.277 33.55 61.44 ;
      END
   END n_80400

   PIN n_80415
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.266 61.277 129.294 61.44 ;
      END
   END n_80415

   PIN n_80418
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.786 61.277 140.814 61.44 ;
      END
   END n_80418

   PIN n_80430
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.37 61.277 144.398 61.44 ;
      END
   END n_80430

   PIN n_80431
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.85 61.277 140.878 61.44 ;
      END
   END n_80431

   PIN n_80488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.138 61.277 33.166 61.44 ;
      END
   END n_80488

   PIN n_80498
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.026 61.277 135.054 61.44 ;
      END
   END n_80498

   PIN n_80510
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.314 0.0 83.342 0.163 ;
      END
   END n_80510

   PIN n_80531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.57 61.277 43.598 61.44 ;
      END
   END n_80531

   PIN n_80539
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.538 61.277 135.566 61.44 ;
      END
   END n_80539

   PIN n_80547
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.722 61.277 44.75 61.44 ;
      END
   END n_80547

   PIN n_80556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.61 61.277 98.638 61.44 ;
      END
   END n_80556

   PIN n_80583
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.274 61.277 36.302 61.44 ;
      END
   END n_80583

   PIN n_80588
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.698 61.277 107.726 61.44 ;
      END
   END n_80588

   PIN n_80590
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.602 61.277 79.63 61.44 ;
      END
   END n_80590

   PIN n_80591
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.394 61.277 89.422 61.44 ;
      END
   END n_80591

   PIN n_80614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.378 0.0 83.406 0.163 ;
      END
   END n_80614

   PIN n_80628
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.65 0.0 81.678 0.163 ;
      END
   END n_80628

   PIN n_80639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.482 61.277 130.51 61.44 ;
      END
   END n_80639

   PIN n_80697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 80.69 61.277 80.718 61.44 ;
      END
   END n_80697

   PIN n_80699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.074 61.277 105.102 61.44 ;
      END
   END n_80699

   PIN n_80702
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.074 61.277 33.102 61.44 ;
      END
   END n_80702

   PIN n_80790
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.114 61.277 32.142 61.44 ;
      END
   END n_80790

   PIN n_80811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.586 61.277 33.614 61.44 ;
      END
   END n_80811

   PIN n_80846
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.522 61.277 57.55 61.44 ;
      END
   END n_80846

   PIN n_80849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.77 61.277 102.798 61.44 ;
      END
   END n_80849

   PIN n_80852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.634 61.277 67.662 61.44 ;
      END
   END n_80852

   PIN n_80863
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.37 61.277 64.398 61.44 ;
      END
   END n_80863

   PIN n_80893
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.498 61.277 56.526 61.44 ;
      END
   END n_80893

   PIN n_81063
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.186 0.163 11.214 ;
      END
   END n_81063

   PIN n_81066
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.25 61.277 99.278 61.44 ;
      END
   END n_81066

   PIN n_81087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.754 61.277 144.782 61.44 ;
      END
   END n_81087

   PIN n_81098
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.338 61.277 52.366 61.44 ;
      END
   END n_81098

   PIN n_81123
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.626 0.163 16.654 ;
      END
   END n_81123

   PIN n_81247
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END n_81247

   PIN n_81358
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.962 0.163 6.99 ;
      END
   END n_81358

   PIN n_81557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.762 0.163 11.79 ;
      END
   END n_81557

   PIN n_81575
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.418 61.277 106.446 61.44 ;
      END
   END n_81575

   PIN n_81588
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.066 61.277 78.094 61.44 ;
      END
   END n_81588

   PIN n_81589
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.002 61.277 78.03 61.44 ;
      END
   END n_81589

   PIN n_81643
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.57 61.277 83.598 61.44 ;
      END
   END n_81643

   PIN n_81647
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.378 61.277 99.406 61.44 ;
      END
   END n_81647

   PIN n_81691
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.466 0.163 12.494 ;
      END
   END n_81691

   PIN n_81748
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.562 61.277 32.59 61.44 ;
      END
   END n_81748

   PIN n_81769
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 73.138 61.277 73.166 61.44 ;
      END
   END n_81769

   PIN n_81897
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.21 0.163 12.238 ;
      END
   END n_81897

   PIN n_81902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.802 61.277 106.83 61.44 ;
      END
   END n_81902

   PIN n_81922
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.418 0.163 26.446 ;
      END
   END n_81922

   PIN n_81929
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.034 0.0 18.062 0.163 ;
      END
   END n_81929

   PIN n_81945
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.666 0.163 7.694 ;
      END
   END n_81945

   PIN n_81985
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.282 61.277 95.31 61.44 ;
      END
   END n_81985

   PIN n_82008
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.906 61.277 105.934 61.44 ;
      END
   END n_82008

   PIN n_82020
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.882 0.163 16.91 ;
      END
   END n_82020

   PIN n_82088
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.282 0.163 15.31 ;
      END
   END n_82088

   PIN n_82097
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.602 61.277 103.63 61.44 ;
      END
   END n_82097

   PIN n_82121
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.858 0.163 7.886 ;
      END
   END n_82121

   PIN n_82123
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.586 61.277 25.614 61.44 ;
      END
   END n_82123

   PIN n_82211
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.218 61.277 95.246 61.44 ;
      END
   END n_82211

   PIN n_82213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.066 61.277 86.094 61.44 ;
      END
   END n_82213

   PIN n_82220
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.058 61.277 91.086 61.44 ;
      END
   END n_82220

   PIN n_82255
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.282 0.163 7.31 ;
      END
   END n_82255

   PIN n_82257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.122 0.163 11.15 ;
      END
   END n_82257

   PIN n_82288
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.29 0.163 2.318 ;
      END
   END n_82288

   PIN n_82318
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.898 61.277 86.926 61.44 ;
      END
   END n_82318

   PIN n_82322
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.802 61.277 90.83 61.44 ;
      END
   END n_82322

   PIN n_82361
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.306 0.163 16.334 ;
      END
   END n_82361

   PIN n_82385
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.962 0.163 14.99 ;
      END
   END n_82385

   PIN n_82411
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.426 61.277 77.454 61.44 ;
      END
   END n_82411

   PIN n_82502
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.218 61.277 87.246 61.44 ;
      END
   END n_82502

   PIN n_82519
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.29 0.163 26.318 ;
      END
   END n_82519

   PIN n_82533
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.57 0.163 35.598 ;
      END
   END n_82533

   PIN n_82546
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.442 61.277 91.47 61.44 ;
      END
   END n_82546

   PIN n_82552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.362 61.277 101.39 61.44 ;
      END
   END n_82552

   PIN n_82605
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.69 0.163 16.718 ;
      END
   END n_82605

   PIN n_82608
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.514 61.277 102.542 61.44 ;
      END
   END n_82608

   PIN n_82617
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.362 61.277 29.39 61.44 ;
      END
   END n_82617

   PIN n_82646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.034 0.163 26.062 ;
      END
   END n_82646

   PIN n_82651
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.338 61.277 20.366 61.44 ;
      END
   END n_82651

   PIN n_82652
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.274 61.277 20.302 61.44 ;
      END
   END n_82652

   PIN n_82657
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.578 0.163 30.606 ;
      END
   END n_82657

   PIN n_82727
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.69 61.277 56.718 61.44 ;
      END
   END n_82727

   PIN n_82772
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.866 0.0 114.894 0.163 ;
      END
   END n_82772

   PIN n_82856
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.082 61.277 60.11 61.44 ;
      END
   END n_82856

   PIN n_82929
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.578 61.277 6.606 61.44 ;
      END
   END n_82929

   PIN n_82932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.89 61.277 67.918 61.44 ;
      END
   END n_82932

   PIN n_82973
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 146.098 61.277 146.126 61.44 ;
      END
   END n_82973

   PIN n_83218
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 144.562 61.277 144.59 61.44 ;
      END
   END n_83218

   PIN n_83282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.794 61.277 71.822 61.44 ;
      END
   END n_83282

   PIN n_83405
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.69 61.277 152.718 61.44 ;
      END
   END n_83405

   PIN n_83632
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 141.042 61.277 141.07 61.44 ;
      END
   END n_83632

   PIN stage2_out_3251
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.594 61.277 20.622 61.44 ;
      END
   END stage2_out_3251

   PIN stage2_out_3285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.602 61.277 71.63 61.44 ;
      END
   END stage2_out_3285

   PIN u1_L14_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.114 61.277 64.142 61.44 ;
      END
   END u1_L14_6_

   PIN u1_L14_reg_29__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.106 61.277 29.134 61.44 ;
      END
   END u1_L14_reg_29__Q

   PIN u2_IP_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.666 61.277 15.694 61.44 ;
      END
   END u2_IP_1_

   PIN u2_IP_64__1283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.522 61.277 25.55 61.44 ;
      END
   END u2_IP_64__1283

   PIN u2_IP_64__1287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.026 61.277 31.054 61.44 ;
      END
   END u2_IP_64__1287

   PIN u2_IP_64__1290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.01 61.277 41.038 61.44 ;
      END
   END u2_IP_64__1290

   PIN u2_L0_21_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.97 61.277 113.998 61.44 ;
      END
   END u2_L0_21_

   PIN u2_L0_22_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.762 61.277 11.79 61.44 ;
      END
   END u2_L0_22_

   PIN u2_L12_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 118.962 61.277 118.99 61.44 ;
      END
   END u2_L12_15_

   PIN u2_L12_21_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.73 61.277 111.758 61.44 ;
      END
   END u2_L12_21_

   PIN u2_L12_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.194 61.277 110.222 61.44 ;
      END
   END u2_L12_5_

   PIN u2_L13_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.346 0.163 15.374 ;
      END
   END u2_L13_23_

   PIN u2_L13_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.658 0.0 44.686 0.163 ;
      END
   END u2_L13_28_

   PIN u2_L1_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.898 61.277 30.926 61.44 ;
      END
   END u2_L1_14_

   PIN u2_L1_25_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.202 61.277 33.23 61.44 ;
      END
   END u2_L1_25_

   PIN u2_L2_reg_7__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.474 61.277 71.502 61.44 ;
      END
   END u2_L2_reg_7__Q

   PIN u2_R0_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.562 61.277 48.59 61.44 ;
      END
   END u2_R0_28_

   PIN u2_R0_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.666 61.277 23.694 61.44 ;
      END
   END u2_R0_8_

   PIN u2_R11_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.634 61.277 75.662 61.44 ;
      END
   END u2_R11_5_

   PIN u2_R12_31_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.85 61.277 44.878 61.44 ;
      END
   END u2_R12_31_

   PIN u2_R13_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 156.466 61.277 156.494 61.44 ;
      END
   END u2_R13_15_

   PIN u2_R13_27_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.81 61.277 117.838 61.44 ;
      END
   END u2_R13_27_

   PIN u2_R14_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 156.21 61.277 156.238 61.44 ;
      END
   END u2_R14_6_

   PIN u2_R1_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.514 61.277 62.542 61.44 ;
      END
   END u2_R1_12_

   PIN u2_R1_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.314 61.277 75.342 61.44 ;
      END
   END u2_R1_7_

   PIN u2_R2_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.754 61.277 40.782 61.44 ;
      END
   END u2_R2_14_

   PIN u2_R2_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.258 61.277 14.286 61.44 ;
      END
   END u2_R2_23_

   PIN u2_R2_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.506 61.277 75.534 61.44 ;
      END
   END u2_R2_28_

   PIN u2_R3_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.802 0.0 90.83 0.163 ;
      END
   END u2_R3_11_

   PIN u2_R3_18_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.658 0.0 124.686 0.163 ;
      END
   END u2_R3_18_

   PIN u2_desIn_r_reg_12__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.77 61.277 22.798 61.44 ;
      END
   END u2_desIn_r_reg_12__Q

   PIN u2_key_r_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.274 61.277 52.302 61.44 ;
      END
   END u2_key_r_14_

   PIN u2_key_r_30_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.21 61.277 52.238 61.44 ;
      END
   END u2_key_r_30_

   PIN u2_key_r_43_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.698 61.277 67.726 61.44 ;
      END
   END u2_key_r_43_

   PIN u2_uk_K_r_222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.722 61.277 44.75 61.44 ;
      END
   END u2_uk_K_r_222

   PIN u2_uk_K_r_365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.49 61.277 29.518 61.44 ;
      END
   END u2_uk_K_r_365

   PIN u2_uk_K_r_380
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.818 61.277 64.846 61.44 ;
      END
   END u2_uk_K_r_380

   PIN u2_uk_K_r_420
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.826 61.277 75.854 61.44 ;
      END
   END u2_uk_K_r_420

   PIN FE_OFN1065_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.658 61.358 52.686 61.44 ;
      END
   END FE_OFN1065_n_116

   PIN FE_OFN1078_n_80338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.226 61.277 138.254 61.44 ;
      END
   END FE_OFN1078_n_80338

   PIN FE_OFN1107_n_20850
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.634 61.277 67.662 61.44 ;
      END
   END FE_OFN1107_n_20850

   PIN FE_OFN1113_n_21429
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.634 61.277 51.662 61.44 ;
      END
   END FE_OFN1113_n_21429

   PIN FE_OFN1151_n_14527
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.21 61.277 60.238 61.44 ;
      END
   END FE_OFN1151_n_14527

   PIN FE_OFN1237_n_19800
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.418 0.0 106.446 0.163 ;
      END
   END FE_OFN1237_n_19800

   PIN FE_OFN1313_n_108168
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 143.154 61.358 143.182 61.44 ;
      END
   END FE_OFN1313_n_108168

   PIN FE_OFN1328_n_82601
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.442 0.163 35.47 ;
      END
   END FE_OFN1328_n_82601

   PIN FE_OFN15_n_106405
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.674 0.0 98.702 0.163 ;
      END
   END FE_OFN15_n_106405

   PIN FE_OFN1820_n_13272
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.394 61.277 25.422 61.44 ;
      END
   END FE_OFN1820_n_13272

   PIN FE_OFN1913_n_78988
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.21 61.277 52.238 61.44 ;
      END
   END FE_OFN1913_n_78988

   PIN FE_OFN217_n_15153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.938 61.277 69.966 61.44 ;
      END
   END FE_OFN217_n_15153

   PIN FE_OFN2233_n_75724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.29 61.277 18.318 61.44 ;
      END
   END FE_OFN2233_n_75724

   PIN FE_OFN2249_n_82961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.17 61.277 77.198 61.44 ;
      END
   END FE_OFN2249_n_82961

   PIN FE_OFN2252_n_80982
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.274 61.277 60.302 61.44 ;
      END
   END FE_OFN2252_n_80982

   PIN FE_OFN244_n_79557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.146 61.277 60.174 61.44 ;
      END
   END FE_OFN244_n_79557

   PIN FE_OFN249_n_79888
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.074 61.277 33.102 61.44 ;
      END
   END FE_OFN249_n_79888

   PIN FE_OFN2516_n_15149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.738 61.277 98.766 61.44 ;
      END
   END FE_OFN2516_n_15149

   PIN FE_OFN255_n_80260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.058 61.277 91.086 61.44 ;
      END
   END FE_OFN255_n_80260

   PIN FE_OFN257_n_79862
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.898 61.277 86.926 61.44 ;
      END
   END FE_OFN257_n_79862

   PIN FE_OFN273_n_75824
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.162 61.277 18.19 61.44 ;
      END
   END FE_OFN273_n_75824

   PIN FE_OFN2762_n_107068
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 144.69 61.277 144.718 61.44 ;
      END
   END FE_OFN2762_n_107068

   PIN FE_OFN2801_n_104989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.834 0.163 30.862 ;
      END
   END FE_OFN2801_n_104989

   PIN FE_OFN2803_n_118632
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.498 61.358 120.526 61.44 ;
      END
   END FE_OFN2803_n_118632

   PIN FE_OFN3160_n_104975
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.69 61.277 8.718 61.44 ;
      END
   END FE_OFN3160_n_104975

   PIN FE_OFN3253_n_39
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.53 61.358 52.558 61.44 ;
      END
   END FE_OFN3253_n_39

   PIN FE_OFN3491_n_83012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.402 61.277 68.43 61.44 ;
      END
   END FE_OFN3491_n_83012

   PIN FE_OFN3495_n_75992
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.562 61.277 48.59 61.44 ;
      END
   END FE_OFN3495_n_75992

   PIN FE_OFN3544_n_105148
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.562 61.277 40.59 61.44 ;
      END
   END FE_OFN3544_n_105148

   PIN FE_OFN3551_n_81000
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.378 61.277 59.406 61.44 ;
      END
   END FE_OFN3551_n_81000

   PIN FE_OFN3553_n_108480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.786 61.277 156.814 61.44 ;
      END
   END FE_OFN3553_n_108480

   PIN FE_OFN4399_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.154 61.358 31.182 61.44 ;
      END
   END FE_OFN4399_decrypt

   PIN FE_OFN4400_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.362 61.358 69.39 61.44 ;
      END
   END FE_OFN4400_decrypt

   PIN FE_OFN821_n_20858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.09 61.277 39.118 61.44 ;
      END
   END FE_OFN821_n_20858

   PIN FE_OFN865_n_15132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.954 61.277 99.982 61.44 ;
      END
   END FE_OFN865_n_15132

   PIN g191933_p1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 22.386 0.163 22.414 ;
      END
   END g191933_p1

   PIN g192018_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 165.746 61.277 165.774 61.44 ;
      END
   END g192018_da

   PIN g192018_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 165.81 61.277 165.838 61.44 ;
      END
   END g192018_db

   PIN g193190_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.298 61.277 125.326 61.44 ;
      END
   END g193190_p

   PIN g194055_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 144.626 61.277 144.654 61.44 ;
      END
   END g194055_da

   PIN g194055_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.626 61.277 144.654 61.44 ;
      END
   END g194055_db

   PIN g194626_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.794 61.277 79.822 61.44 ;
      END
   END g194626_p

   PIN g197833_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.194 0.0 110.222 0.163 ;
      END
   END g197833_da

   PIN g198664_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.69 61.277 72.718 61.44 ;
      END
   END g198664_p

   PIN g215918_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.746 61.277 69.774 61.44 ;
      END
   END g215918_p

   PIN g216302_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.978 61.277 69.006 61.44 ;
      END
   END g216302_db

   PIN g216302_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.538 61.277 63.566 61.44 ;
      END
   END g216302_sb

   PIN g216515_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.162 61.277 98.19 61.44 ;
      END
   END g216515_da

   PIN g216515_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.226 61.277 98.254 61.44 ;
      END
   END g216515_db

   PIN g216746_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.282 61.277 79.31 61.44 ;
      END
   END g216746_sb

   PIN g217136_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.602 61.277 23.63 61.44 ;
      END
   END g217136_p

   PIN g217299_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.314 61.277 83.342 61.44 ;
      END
   END g217299_p

   PIN g218012_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.194 0.0 14.222 0.163 ;
      END
   END g218012_p

   PIN g219309_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.69 61.277 40.718 61.44 ;
      END
   END g219309_p

   PIN g219396_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.642 61.277 94.67 61.44 ;
      END
   END g219396_p

   PIN g219482_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.33 61.277 33.358 61.44 ;
      END
   END g219482_p

   PIN g219847_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.946 61.277 40.974 61.44 ;
      END
   END g219847_p

   PIN g220720_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.29 61.277 114.318 61.44 ;
      END
   END g220720_da

   PIN g220720_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.458 61.277 25.486 61.44 ;
      END
   END g220720_db

   PIN g220874_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.706 61.277 22.734 61.44 ;
      END
   END g220874_db

   PIN g220874_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.21 61.277 20.238 61.44 ;
      END
   END g220874_sb

   PIN g222231_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.162 61.277 18.19 61.44 ;
      END
   END g222231_p

   PIN g222770_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.618 61.277 21.646 61.44 ;
      END
   END g222770_db

   PIN g222770_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.562 61.277 16.59 61.44 ;
      END
   END g222770_sb

   PIN g223067_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.97 61.277 25.998 61.44 ;
      END
   END g223067_da

   PIN g223067_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.034 61.277 26.062 61.44 ;
      END
   END g223067_db

   PIN g223067_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.65 61.277 25.678 61.44 ;
      END
   END g223067_sb

   PIN g223077_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.186 61.277 35.214 61.44 ;
      END
   END g223077_db

   PIN g223077_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.106 61.277 37.134 61.44 ;
      END
   END g223077_sb

   PIN g224248_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.178 61.277 16.206 61.44 ;
      END
   END g224248_db

   PIN g288145_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.242 61.277 56.27 61.44 ;
      END
   END g288145_p

   PIN g288651_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.314 61.277 27.342 61.44 ;
      END
   END g288651_p

   PIN g322456_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.978 61.277 45.006 61.44 ;
      END
   END g322456_sb

   PIN g322683_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.882 61.277 144.91 61.44 ;
      END
   END g322683_da

   PIN g322683_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.818 61.277 144.846 61.44 ;
      END
   END g322683_db

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.202 61.277 41.23 61.44 ;
      END
   END ispd_clk

   PIN key_c_r_30__2103
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.706 61.277 70.734 61.44 ;
      END
   END key_c_r_30__2103

   PIN key_c_r_32__2208
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.226 0.0 90.254 0.163 ;
      END
   END key_c_r_32__2208

   PIN key_c_r_32__2214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.57 61.277 75.598 61.44 ;
      END
   END key_c_r_32__2214

   PIN key_c_r_32__2243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.346 61.277 79.374 61.44 ;
      END
   END key_c_r_32__2243

   PIN key_c_r_33__30_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.466 0.163 44.494 ;
      END
   END key_c_r_33__30_

   PIN n_100299
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.738 61.277 74.766 61.44 ;
      END
   END n_100299

   PIN n_100477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.546 61.277 90.574 61.44 ;
      END
   END n_100477

   PIN n_100495
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.994 61.277 83.022 61.44 ;
      END
   END n_100495

   PIN n_100662
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.17 61.277 77.198 61.44 ;
      END
   END n_100662

   PIN n_100714
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.314 61.277 83.342 61.44 ;
      END
   END n_100714

   PIN n_100761
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.354 61.277 90.382 61.44 ;
      END
   END n_100761

   PIN n_100762
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.162 61.277 90.19 61.44 ;
      END
   END n_100762

   PIN n_101445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 125.042 61.277 125.07 61.44 ;
      END
   END n_101445

   PIN n_101500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 136.946 61.277 136.974 61.44 ;
      END
   END n_101500

   PIN n_101504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.882 61.277 128.91 61.44 ;
      END
   END n_101504

   PIN n_101636
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 125.106 61.277 125.134 61.44 ;
      END
   END n_101636

   PIN n_101645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 131.378 61.277 131.406 61.44 ;
      END
   END n_101645

   PIN n_101699
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 140.786 61.277 140.814 61.44 ;
      END
   END n_101699

   PIN n_101768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 128.178 61.277 128.206 61.44 ;
      END
   END n_101768

   PIN n_101913
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 122.546 61.277 122.574 61.44 ;
      END
   END n_101913

   PIN n_102201
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 140.914 61.277 140.942 61.44 ;
      END
   END n_102201

   PIN n_102880
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 156.338 61.277 156.366 61.44 ;
      END
   END n_102880

   PIN n_102908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.922 61.277 63.95 61.44 ;
      END
   END n_102908

   PIN n_102997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.602 61.277 79.63 61.44 ;
      END
   END n_102997

   PIN n_103008
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.85 0.0 44.878 0.163 ;
      END
   END n_103008

   PIN n_103115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.754 61.277 48.782 61.44 ;
      END
   END n_103115

   PIN n_103266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.994 61.277 91.022 61.44 ;
      END
   END n_103266

   PIN n_103664
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.482 61.277 90.51 61.44 ;
      END
   END n_103664

   PIN n_103670
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.25 61.277 83.278 61.44 ;
      END
   END n_103670

   PIN n_103671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.834 61.277 86.862 61.44 ;
      END
   END n_103671

   PIN n_103694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.986 61.277 88.014 61.44 ;
      END
   END n_103694

   PIN n_103802
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.778 61.277 81.806 61.44 ;
      END
   END n_103802

   PIN n_103837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.77 61.277 86.798 61.44 ;
      END
   END n_103837

   PIN n_103855
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.162 61.277 90.19 61.44 ;
      END
   END n_103855

   PIN n_103882
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.202 61.277 81.23 61.44 ;
      END
   END n_103882

   PIN n_103972
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.994 61.277 83.022 61.44 ;
      END
   END n_103972

   PIN n_103998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.706 61.277 86.734 61.44 ;
      END
   END n_103998

   PIN n_104090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.106 61.277 85.134 61.44 ;
      END
   END n_104090

   PIN n_104111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.362 61.277 85.39 61.44 ;
      END
   END n_104111

   PIN n_104147
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.482 61.277 90.51 61.44 ;
      END
   END n_104147

   PIN n_104148
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.45 61.277 78.478 61.44 ;
      END
   END n_104148

   PIN n_104284
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.642 61.277 86.67 61.44 ;
      END
   END n_104284

   PIN n_104373
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.186 61.277 83.214 61.44 ;
      END
   END n_104373

   PIN n_104411
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.578 61.277 86.606 61.44 ;
      END
   END n_104411

   PIN n_104493
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.618 61.277 85.646 61.44 ;
      END
   END n_104493

   PIN n_104505
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.65 61.277 81.678 61.44 ;
      END
   END n_104505

   PIN n_104520
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.122 61.277 83.15 61.44 ;
      END
   END n_104520

   PIN n_104588
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.17 61.277 85.198 61.44 ;
      END
   END n_104588

   PIN n_104625
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.386 61.277 78.414 61.44 ;
      END
   END n_104625

   PIN n_104873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.402 61.277 148.43 61.44 ;
      END
   END n_104873

   PIN n_105003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.074 61.277 73.102 61.44 ;
      END
   END n_105003

   PIN n_105099
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.93 61.277 82.958 61.44 ;
      END
   END n_105099

   PIN n_105150
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.162 61.277 114.19 61.44 ;
      END
   END n_105150

   PIN n_105176
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.122 0.163 19.15 ;
      END
   END n_105176

   PIN n_105284
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.058 0.163 19.086 ;
      END
   END n_105284

   PIN n_105286
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.738 0.163 26.766 ;
      END
   END n_105286

   PIN n_105287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.706 0.082 30.734 ;
      END
   END n_105287

   PIN n_105353
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.442 0.163 19.47 ;
      END
   END n_105353

   PIN n_105423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.794 0.0 71.822 0.163 ;
      END
   END n_105423

   PIN n_105424
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.17 61.277 69.198 61.44 ;
      END
   END n_105424

   PIN n_105451
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.746 0.163 21.774 ;
      END
   END n_105451

   PIN n_105486
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.338 61.277 116.366 61.44 ;
      END
   END n_105486

   PIN n_105503
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.082 0.0 68.11 0.163 ;
      END
   END n_105503

   PIN n_105531
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.938 0.163 21.966 ;
      END
   END n_105531

   PIN n_105540
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.826 0.0 67.854 0.163 ;
      END
   END n_105540

   PIN n_105541
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.834 0.0 70.862 0.163 ;
      END
   END n_105541

   PIN n_105547
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.674 0.163 26.702 ;
      END
   END n_105547

   PIN n_105552
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.778 61.277 161.806 61.44 ;
      END
   END n_105552

   PIN n_105593
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.554 0.0 61.582 0.163 ;
      END
   END n_105593

   PIN n_105596
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.994 0.0 91.022 0.163 ;
      END
   END n_105596

   PIN n_105632
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.762 0.0 67.79 0.163 ;
      END
   END n_105632

   PIN n_105634
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.25 0.163 19.278 ;
      END
   END n_105634

   PIN n_105645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.346 0.0 63.374 0.163 ;
      END
   END n_105645

   PIN n_105648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.426 61.277 117.454 61.44 ;
      END
   END n_105648

   PIN n_105678
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.714 61.277 161.742 61.44 ;
      END
   END n_105678

   PIN n_105694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.906 0.163 25.934 ;
      END
   END n_105694

   PIN n_105696
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.074 0.0 73.102 0.163 ;
      END
   END n_105696

   PIN n_105707
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.466 61.277 116.494 61.44 ;
      END
   END n_105707

   PIN n_105715
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.986 0.0 80.014 0.163 ;
      END
   END n_105715

   PIN n_105739
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.242 0.0 64.27 0.163 ;
      END
   END n_105739

   PIN n_105749
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.474 0.0 79.502 0.163 ;
      END
   END n_105749

   PIN n_105788
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.322 0.163 30.35 ;
      END
   END n_105788

   PIN n_105875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.682 0.163 21.71 ;
      END
   END n_105875

   PIN n_105910
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.45 0.163 22.478 ;
      END
   END n_105910

   PIN n_105912
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.85 0.0 68.878 0.163 ;
      END
   END n_105912

   PIN n_105916
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.73 0.0 71.758 0.163 ;
      END
   END n_105916

   PIN n_105937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.618 0.163 21.646 ;
      END
   END n_105937

   PIN n_105995
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.698 0.0 75.726 0.163 ;
      END
   END n_105995

   PIN n_106012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.618 61.277 125.646 61.44 ;
      END
   END n_106012

   PIN n_106014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.306 61.277 120.334 61.44 ;
      END
   END n_106014

   PIN n_106037
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.098 0.163 26.126 ;
      END
   END n_106037

   PIN n_106057
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.426 61.277 125.454 61.44 ;
      END
   END n_106057

   PIN n_106089
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.554 0.163 21.582 ;
      END
   END n_106089

   PIN n_106090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.994 0.163 19.022 ;
      END
   END n_106090

   PIN n_106099
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.61 0.163 26.638 ;
      END
   END n_106099

   PIN n_106148
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.978 61.277 117.006 61.44 ;
      END
   END n_106148

   PIN n_106153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.93 0.163 18.958 ;
      END
   END n_106153

   PIN n_106158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.434 0.0 56.462 0.163 ;
      END
   END n_106158

   PIN n_106159
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.594 0.0 52.622 0.163 ;
      END
   END n_106159

   PIN n_106162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.642 0.163 22.67 ;
      END
   END n_106162

   PIN n_106163
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.49 0.163 21.518 ;
      END
   END n_106163

   PIN n_106166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.578 0.163 22.606 ;
      END
   END n_106166

   PIN n_106171
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.186 0.0 59.214 0.163 ;
      END
   END n_106171

   PIN n_106182
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.058 61.277 123.086 61.44 ;
      END
   END n_106182

   PIN n_106184
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 160.818 61.277 160.846 61.44 ;
      END
   END n_106184

   PIN n_106194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.082 0.0 60.11 0.163 ;
      END
   END n_106194

   PIN n_106196
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.498 0.163 16.526 ;
      END
   END n_106196

   PIN n_106200
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.954 0.0 67.982 0.163 ;
      END
   END n_106200

   PIN n_106207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.538 61.277 127.566 61.44 ;
      END
   END n_106207

   PIN n_106208
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.522 61.277 121.55 61.44 ;
      END
   END n_106208

   PIN n_106220
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.866 0.163 18.894 ;
      END
   END n_106220

   PIN n_106224
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.69 0.0 48.718 0.163 ;
      END
   END n_106224

   PIN n_106247
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.93 61.277 122.958 61.44 ;
      END
   END n_106247

   PIN n_106253
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.378 0.163 19.406 ;
      END
   END n_106253

   PIN n_106258
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.514 0.163 22.542 ;
      END
   END n_106258

   PIN n_106273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.314 0.163 19.342 ;
      END
   END n_106273

   PIN n_106306
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.234 61.277 125.262 61.44 ;
      END
   END n_106306

   PIN n_106327
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.834 0.163 22.862 ;
      END
   END n_106327

   PIN n_106329
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.802 0.163 26.83 ;
      END
   END n_106329

   PIN n_106337
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 19.186 0.163 19.214 ;
      END
   END n_106337

   PIN n_106361
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.434 0.0 64.462 0.163 ;
      END
   END n_106361

   PIN n_106445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.034 0.0 66.062 0.163 ;
      END
   END n_106445

   PIN n_106450
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.922 0.0 63.95 0.163 ;
      END
   END n_106450

   PIN n_106452
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.802 0.163 18.83 ;
      END
   END n_106452

   PIN n_106488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.866 61.277 122.894 61.44 ;
      END
   END n_106488

   PIN n_106510
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.474 61.277 119.502 61.44 ;
      END
   END n_106510

   PIN n_106526
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.426 0.163 21.454 ;
      END
   END n_106526

   PIN n_106531
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.938 0.0 45.966 0.163 ;
      END
   END n_106531

   PIN n_106533
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.554 61.277 125.582 61.44 ;
      END
   END n_106533

   PIN n_106568
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.37 0.0 56.398 0.163 ;
      END
   END n_106568

   PIN n_106586
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.738 0.0 58.766 0.163 ;
      END
   END n_106586

   PIN n_106596
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.218 0.0 87.246 0.163 ;
      END
   END n_106596

   PIN n_106597
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.53 0.0 52.558 0.163 ;
      END
   END n_106597

   PIN n_106601
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.378 0.0 51.406 0.163 ;
      END
   END n_106601

   PIN n_106603
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.226 0.163 2.254 ;
      END
   END n_106603

   PIN n_106608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.858 0.0 63.886 0.163 ;
      END
   END n_106608

   PIN n_106629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.458 61.277 121.486 61.44 ;
      END
   END n_106629

   PIN n_106649
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.738 0.163 18.766 ;
      END
   END n_106649

   PIN n_106661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.538 61.277 119.566 61.44 ;
      END
   END n_106661

   PIN n_106663
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.634 0.0 75.662 0.163 ;
      END
   END n_106663

   PIN n_106710
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.49 61.277 125.518 61.44 ;
      END
   END n_106710

   PIN n_106714
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.402 0.163 12.43 ;
      END
   END n_106714

   PIN n_106751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.394 61.277 121.422 61.44 ;
      END
   END n_106751

   PIN n_106817
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.978 0.0 45.006 0.163 ;
      END
   END n_106817

   PIN n_106818
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.402 61.277 156.43 61.44 ;
      END
   END n_106818

   PIN n_106840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.914 0.0 44.942 0.163 ;
      END
   END n_106840

   PIN n_106900
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 160.306 61.277 160.334 61.44 ;
      END
   END n_106900

   PIN n_107024
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 165.426 61.277 165.454 61.44 ;
      END
   END n_107024

   PIN n_107054
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 16.306 167.36 16.334 ;
      END
   END n_107054

   PIN n_107067
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.698 61.277 155.726 61.44 ;
      END
   END n_107067

   PIN n_107081
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.498 61.277 160.526 61.44 ;
      END
   END n_107081

   PIN n_107097
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.882 61.277 160.91 61.44 ;
      END
   END n_107097

   PIN n_107129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.09 61.277 151.118 61.44 ;
      END
   END n_107129

   PIN n_107136
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.05 61.277 152.078 61.44 ;
      END
   END n_107136

   PIN n_107146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 155.954 61.277 155.982 61.44 ;
      END
   END n_107146

   PIN n_107190
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 149.682 61.358 149.71 61.44 ;
      END
   END n_107190

   PIN n_107250
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 160.37 61.277 160.398 61.44 ;
      END
   END n_107250

   PIN n_107253
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.626 61.277 160.654 61.44 ;
      END
   END n_107253

   PIN n_107341
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.69 61.277 160.718 61.44 ;
      END
   END n_107341

   PIN n_107345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.122 0.0 163.15 0.163 ;
      END
   END n_107345

   PIN n_107369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 45.042 167.36 45.07 ;
      END
   END n_107369

   PIN n_107412
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.754 61.277 160.782 61.44 ;
      END
   END n_107412

   PIN n_107462
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 39.922 167.36 39.95 ;
      END
   END n_107462

   PIN n_107486
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 44.466 167.36 44.494 ;
      END
   END n_107486

   PIN n_107495
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.466 61.277 164.494 61.44 ;
      END
   END n_107495

   PIN n_107519
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 30.386 167.36 30.414 ;
      END
   END n_107519

   PIN n_107577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.978 0.0 141.006 0.163 ;
      END
   END n_107577

   PIN n_107602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.434 61.277 160.462 61.44 ;
      END
   END n_107602

   PIN n_107611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.954 61.277 155.982 61.44 ;
      END
   END n_107611

   PIN n_107634
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.042 0.0 149.07 0.163 ;
      END
   END n_107634

   PIN n_107640
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.818 61.277 160.846 61.44 ;
      END
   END n_107640

   PIN n_107641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 44.402 167.36 44.43 ;
      END
   END n_107641

   PIN n_107652
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 160.242 61.277 160.27 61.44 ;
      END
   END n_107652

   PIN n_107656
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 22.962 167.36 22.99 ;
      END
   END n_107656

   PIN n_107660
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.09 61.277 159.118 61.44 ;
      END
   END n_107660

   PIN n_107674
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 54.002 167.36 54.03 ;
      END
   END n_107674

   PIN n_107677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.278 35.442 167.36 35.47 ;
      END
   END n_107677

   PIN n_107723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.338 61.277 148.366 61.44 ;
      END
   END n_107723

   PIN n_107738
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.89 0.0 163.918 0.163 ;
      END
   END n_107738

   PIN n_107746
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.658 61.277 148.686 61.44 ;
      END
   END n_107746

   PIN n_107782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.018 61.277 156.046 61.44 ;
      END
   END n_107782

   PIN n_107829
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.034 0.0 114.062 0.163 ;
      END
   END n_107829

   PIN n_107928
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.082 61.277 156.11 61.44 ;
      END
   END n_107928

   PIN n_107943
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 7.282 167.36 7.31 ;
      END
   END n_107943

   PIN n_107996
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 26.738 167.36 26.766 ;
      END
   END n_107996

   PIN n_108012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.37 61.277 160.398 61.44 ;
      END
   END n_108012

   PIN n_108045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 11.442 167.36 11.47 ;
      END
   END n_108045

   PIN n_108049
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.938 61.277 157.966 61.44 ;
      END
   END n_108049

   PIN n_108137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.21 61.277 156.238 61.44 ;
      END
   END n_108137

   PIN n_108148
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.394 61.277 153.422 61.44 ;
      END
   END n_108148

   PIN n_108191
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.466 61.277 148.494 61.44 ;
      END
   END n_108191

   PIN n_108245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.274 0.0 156.302 0.163 ;
      END
   END n_108245

   PIN n_108254
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.562 61.277 144.59 61.44 ;
      END
   END n_108254

   PIN n_108278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.546 61.277 154.574 61.44 ;
      END
   END n_108278

   PIN n_108295
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 22.898 167.36 22.926 ;
      END
   END n_108295

   PIN n_108407
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 25.906 167.36 25.934 ;
      END
   END n_108407

   PIN n_108410
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 167.197 30.322 167.36 30.35 ;
      END
   END n_108410

   PIN n_108418
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.53 61.277 148.558 61.44 ;
      END
   END n_108418

   PIN n_108449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.722 61.277 148.75 61.44 ;
      END
   END n_108449

   PIN n_108499
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.746 61.277 157.774 61.44 ;
      END
   END n_108499

   PIN n_109142
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.234 61.277 37.262 61.44 ;
      END
   END n_109142

   PIN n_109209
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.762 61.277 35.79 61.44 ;
      END
   END n_109209

   PIN n_116820
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.242 61.277 128.27 61.44 ;
      END
   END n_116820

   PIN n_117788
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.53 61.277 60.558 61.44 ;
      END
   END n_117788

   PIN n_118032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.402 61.277 164.43 61.44 ;
      END
   END n_118032

   PIN n_118355
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.682 61.277 93.71 61.44 ;
      END
   END n_118355

   PIN n_118357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.05 61.277 88.078 61.44 ;
      END
   END n_118357

   PIN n_118359
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.154 61.277 87.182 61.44 ;
      END
   END n_118359

   PIN n_118364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.898 61.277 94.926 61.44 ;
      END
   END n_118364

   PIN n_118371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.378 61.277 91.406 61.44 ;
      END
   END n_118371

   PIN n_118636
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.362 61.277 125.39 61.44 ;
      END
   END n_118636

   PIN n_118642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.682 61.277 117.71 61.44 ;
      END
   END n_118642

   PIN n_118707
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.674 61.277 98.702 61.44 ;
      END
   END n_118707

   PIN n_126097
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.082 61.277 132.11 61.44 ;
      END
   END n_126097

   PIN n_13376
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.706 61.277 30.734 61.44 ;
      END
   END n_13376

   PIN n_13380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.73 61.277 39.758 61.44 ;
      END
   END n_13380

   PIN n_13382
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.514 61.277 46.542 61.44 ;
      END
   END n_13382

   PIN n_13477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.658 61.277 44.686 61.44 ;
      END
   END n_13477

   PIN n_13479
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.658 61.277 44.686 61.44 ;
      END
   END n_13479

   PIN n_13482
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.594 61.277 44.622 61.44 ;
      END
   END n_13482

   PIN n_13488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.994 61.277 35.022 61.44 ;
      END
   END n_13488

   PIN n_13521
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.946 61.277 0.974 61.44 ;
      END
   END n_13521

   PIN n_13606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.69 61.277 40.718 61.44 ;
      END
   END n_13606

   PIN n_13710
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.682 61.277 69.71 61.44 ;
      END
   END n_13710

   PIN n_137147
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.274 0.163 12.302 ;
      END
   END n_137147

   PIN n_137154
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.578 61.277 6.606 61.44 ;
      END
   END n_137154

   PIN n_13741
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.042 61.277 37.07 61.44 ;
      END
   END n_13741

   PIN n_13754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.25 61.277 35.278 61.44 ;
      END
   END n_13754

   PIN n_13841
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.33 61.277 65.358 61.44 ;
      END
   END n_13841

   PIN n_13861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.01 61.277 41.038 61.44 ;
      END
   END n_13861

   PIN n_13872
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.026 61.277 71.054 61.44 ;
      END
   END n_13872

   PIN n_13981
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.818 61.277 56.846 61.44 ;
      END
   END n_13981

   PIN n_14011
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.442 61.277 59.47 61.44 ;
      END
   END n_14011

   PIN n_14014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.626 61.277 56.654 61.44 ;
      END
   END n_14014

   PIN n_14026
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.498 61.277 48.526 61.44 ;
      END
   END n_14026

   PIN n_14129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.29 61.277 42.318 61.44 ;
      END
   END n_14129

   PIN n_14373
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.754 61.277 40.782 61.44 ;
      END
   END n_14373

   PIN n_14379
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.242 61.277 48.27 61.44 ;
      END
   END n_14379

   PIN n_14517
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.458 61.277 57.486 61.44 ;
      END
   END n_14517

   PIN n_14520
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.89 61.277 51.918 61.44 ;
      END
   END n_14520

   PIN n_14525
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.298 61.277 53.326 61.44 ;
      END
   END n_14525

   PIN n_15151
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.594 61.277 52.622 61.44 ;
      END
   END n_15151

   PIN n_15369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.826 61.277 67.854 61.44 ;
      END
   END n_15369

   PIN n_212521
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.25 61.277 51.278 61.44 ;
      END
   END n_212521

   PIN n_21351
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.354 61.277 18.382 61.44 ;
      END
   END n_21351

   PIN n_21398
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.338 61.277 60.366 61.44 ;
      END
   END n_21398

   PIN n_21430
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.722 61.277 52.75 61.44 ;
      END
   END n_21430

   PIN n_75475
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.186 61.277 27.214 61.44 ;
      END
   END n_75475

   PIN n_75713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.962 61.277 30.99 61.44 ;
      END
   END n_75713

   PIN n_75715
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.25 61.277 27.278 61.44 ;
      END
   END n_75715

   PIN n_75770
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.49 61.277 61.518 61.44 ;
      END
   END n_75770

   PIN n_75788
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.074 61.277 49.102 61.44 ;
      END
   END n_75788

   PIN n_76012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.042 61.277 5.07 61.44 ;
      END
   END n_76012

   PIN n_76214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.33 61.358 9.358 61.44 ;
      END
   END n_76214

   PIN n_76298
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.194 61.277 14.222 61.44 ;
      END
   END n_76298

   PIN n_76529
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.49 61.277 21.518 61.44 ;
      END
   END n_76529

   PIN n_76816
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.386 61.277 14.414 61.44 ;
      END
   END n_76816

   PIN n_76865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.186 61.277 3.214 61.44 ;
      END
   END n_76865

   PIN n_76896
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.546 61.277 18.574 61.44 ;
      END
   END n_76896

   PIN n_76931
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.226 61.277 18.254 61.44 ;
      END
   END n_76931

   PIN n_76932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.01 61.277 17.038 61.44 ;
      END
   END n_76932

   PIN n_76935
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.554 61.277 21.582 61.44 ;
      END
   END n_76935

   PIN n_77062
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.074 61.277 17.102 61.44 ;
      END
   END n_77062

   PIN n_77148
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.002 61.277 14.03 61.44 ;
      END
   END n_77148

   PIN n_77280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.41 61.277 7.438 61.44 ;
      END
   END n_77280

   PIN n_77331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.482 61.277 18.51 61.44 ;
      END
   END n_77331

   PIN n_77392
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.066 61.358 14.094 61.44 ;
      END
   END n_77392

   PIN n_77415
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.01 61.277 1.038 61.44 ;
      END
   END n_77415

   PIN n_77416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.194 61.277 14.222 61.44 ;
      END
   END n_77416

   PIN n_77722
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.162 61.277 10.19 61.44 ;
      END
   END n_77722

   PIN n_77723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.914 61.277 12.942 61.44 ;
      END
   END n_77723

   PIN n_77759
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.258 61.277 14.286 61.44 ;
      END
   END n_77759

   PIN n_77771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.066 61.277 14.094 61.44 ;
      END
   END n_77771

   PIN n_77821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.29 61.277 10.318 61.44 ;
      END
   END n_77821

   PIN n_77947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.106 61.277 5.134 61.44 ;
      END
   END n_77947

   PIN n_78815
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.642 61.277 6.67 61.44 ;
      END
   END n_78815

   PIN n_78831
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.466 61.277 52.494 61.44 ;
      END
   END n_78831

   PIN n_78876
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.026 61.277 95.054 61.44 ;
      END
   END n_78876

   PIN n_78916
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.602 61.277 71.63 61.44 ;
      END
   END n_78916

   PIN n_78927
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.978 61.277 37.006 61.44 ;
      END
   END n_78927

   PIN n_78965
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.258 61.277 54.286 61.44 ;
      END
   END n_78965

   PIN n_78977
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.25 61.277 91.278 61.44 ;
      END
   END n_78977

   PIN n_78990
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.754 61.277 56.782 61.44 ;
      END
   END n_78990

   PIN n_78998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.402 61.277 52.43 61.44 ;
      END
   END n_78998

   PIN n_79103
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.314 61.277 51.342 61.44 ;
      END
   END n_79103

   PIN n_79120
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.074 61.277 41.102 61.44 ;
      END
   END n_79120

   PIN n_79137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.186 61.277 91.214 61.44 ;
      END
   END n_79137

   PIN n_79146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.402 61.277 60.43 61.44 ;
      END
   END n_79146

   PIN n_79180
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.258 61.277 110.286 61.44 ;
      END
   END n_79180

   PIN n_79289
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.05 61.277 136.078 61.44 ;
      END
   END n_79289

   PIN n_79305
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.882 61.277 40.91 61.44 ;
      END
   END n_79305

   PIN n_79354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.73 61.277 71.758 61.44 ;
      END
   END n_79354

   PIN n_79364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.026 61.277 87.054 61.44 ;
      END
   END n_79364

   PIN n_79384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.666 61.277 103.694 61.44 ;
      END
   END n_79384

   PIN n_79386
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.066 61.277 46.094 61.44 ;
      END
   END n_79386

   PIN n_79389
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.866 61.277 58.894 61.44 ;
      END
   END n_79389

   PIN n_79393
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.53 61.277 28.558 61.44 ;
      END
   END n_79393

   PIN n_79422
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.978 61.277 93.006 61.44 ;
      END
   END n_79422

   PIN n_79423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.146 61.277 76.174 61.44 ;
      END
   END n_79423

   PIN n_79461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.29 61.277 138.318 61.44 ;
      END
   END n_79461

   PIN n_79469
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.162 61.277 50.19 61.44 ;
      END
   END n_79469

   PIN n_79525
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.314 61.277 91.342 61.44 ;
      END
   END n_79525

   PIN n_79565
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.794 0.0 111.822 0.163 ;
      END
   END n_79565

   PIN n_79566
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.962 61.277 86.99 61.44 ;
      END
   END n_79566

   PIN n_79570
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.658 61.277 28.686 61.44 ;
      END
   END n_79570

   PIN n_79571
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.498 61.277 40.526 61.44 ;
      END
   END n_79571

   PIN n_79575
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.33 61.277 129.358 61.44 ;
      END
   END n_79575

   PIN n_79576
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.074 61.277 41.102 61.44 ;
      END
   END n_79576

   PIN n_79622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.09 61.277 87.118 61.44 ;
      END
   END n_79622

   PIN n_79636
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.474 61.277 79.502 61.44 ;
      END
   END n_79636

   PIN n_79679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.41 61.277 79.438 61.44 ;
      END
   END n_79679

   PIN n_79720
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.794 61.277 103.822 61.44 ;
      END
   END n_79720

   PIN n_79734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.802 61.277 90.83 61.44 ;
      END
   END n_79734

   PIN n_79739
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.93 61.277 90.958 61.44 ;
      END
   END n_79739

   PIN n_79776
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.698 61.277 139.726 61.44 ;
      END
   END n_79776

   PIN n_79781
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.498 61.277 128.526 61.44 ;
      END
   END n_79781

   PIN n_79802
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.89 61.277 75.918 61.44 ;
      END
   END n_79802

   PIN n_79857
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.65 61.277 33.678 61.44 ;
      END
   END n_79857

   PIN n_79870
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.394 61.277 33.422 61.44 ;
      END
   END n_79870

   PIN n_79886
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.682 61.277 37.71 61.44 ;
      END
   END n_79886

   PIN n_79924
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.914 61.277 132.942 61.44 ;
      END
   END n_79924

   PIN n_79933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.33 61.277 137.358 61.44 ;
      END
   END n_79933

   PIN n_79945
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.626 61.277 96.654 61.44 ;
      END
   END n_79945

   PIN n_79963
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.09 61.277 79.118 61.44 ;
      END
   END n_79963

   PIN n_79967
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.298 61.277 37.326 61.44 ;
      END
   END n_79967

   PIN n_80003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.322 61.277 110.35 61.44 ;
      END
   END n_80003

   PIN n_80022
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.698 61.277 43.726 61.44 ;
      END
   END n_80022

   PIN n_80032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.762 61.277 67.79 61.44 ;
      END
   END n_80032

   PIN n_80060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.642 61.277 142.67 61.44 ;
      END
   END n_80060

   PIN n_80067
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.362 61.277 133.39 61.44 ;
      END
   END n_80067

   PIN n_80068
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.682 61.277 133.71 61.44 ;
      END
   END n_80068

   PIN n_80096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.794 61.277 135.822 61.44 ;
      END
   END n_80096

   PIN n_80115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.866 61.277 90.894 61.44 ;
      END
   END n_80115

   PIN n_80137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.018 61.277 108.046 61.44 ;
      END
   END n_80137

   PIN n_80149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.954 61.277 67.982 61.44 ;
      END
   END n_80149

   PIN n_80206
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 130.546 61.358 130.574 61.44 ;
      END
   END n_80206

   PIN n_80245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.85 61.277 132.878 61.44 ;
      END
   END n_80245

   PIN n_80249
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.946 61.277 40.974 61.44 ;
      END
   END n_80249

   PIN n_80253
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.042 61.277 45.07 61.44 ;
      END
   END n_80253

   PIN n_80274
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 140.85 61.277 140.878 61.44 ;
      END
   END n_80274

   PIN n_80282
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.826 61.277 67.854 61.44 ;
      END
   END n_80282

   PIN n_80325
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.69 61.277 136.718 61.44 ;
      END
   END n_80325

   PIN n_80329
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.298 61.277 133.326 61.44 ;
      END
   END n_80329

   PIN n_80387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.866 61.277 90.894 61.44 ;
      END
   END n_80387

   PIN n_80393
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 84.914 61.277 84.942 61.44 ;
      END
   END n_80393

   PIN n_80399
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.466 61.277 100.494 61.44 ;
      END
   END n_80399

   PIN n_80401
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.618 61.277 45.646 61.44 ;
      END
   END n_80401

   PIN n_80404
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.458 61.277 33.486 61.44 ;
      END
   END n_80404

   PIN n_80408
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.138 61.277 129.166 61.44 ;
      END
   END n_80408

   PIN n_80412
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.234 61.277 133.262 61.44 ;
      END
   END n_80412

   PIN n_80425
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.338 61.277 84.366 61.44 ;
      END
   END n_80425

   PIN n_80429
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.818 61.277 136.846 61.44 ;
      END
   END n_80429

   PIN n_80504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.218 61.277 71.246 61.44 ;
      END
   END n_80504

   PIN n_80520
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.362 61.277 37.39 61.44 ;
      END
   END n_80520

   PIN n_80538
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.73 61.277 135.758 61.44 ;
      END
   END n_80538

   PIN n_80551
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.242 61.277 64.27 61.44 ;
      END
   END n_80551

   PIN n_80557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.634 61.277 59.662 61.44 ;
      END
   END n_80557

   PIN n_80619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.394 61.277 25.422 61.44 ;
      END
   END n_80619

   PIN n_80631
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.714 61.277 89.742 61.44 ;
      END
   END n_80631

   PIN n_80640
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.61 61.277 130.638 61.44 ;
      END
   END n_80640

   PIN n_80682
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.122 61.277 99.15 61.44 ;
      END
   END n_80682

   PIN n_80694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.306 61.277 56.334 61.44 ;
      END
   END n_80694

   PIN n_80734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.106 61.277 45.134 61.44 ;
      END
   END n_80734

   PIN n_80743
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.29 61.277 90.318 61.44 ;
      END
   END n_80743

   PIN n_80759
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.906 61.277 49.934 61.44 ;
      END
   END n_80759

   PIN n_80763
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.33 61.277 73.358 61.44 ;
      END
   END n_80763

   PIN n_80777
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.322 61.277 134.35 61.44 ;
      END
   END n_80777

   PIN n_80788
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.25 0.0 83.278 0.163 ;
      END
   END n_80788

   PIN n_80817
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.226 61.277 114.254 61.44 ;
      END
   END n_80817

   PIN n_80905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.37 61.277 56.398 61.44 ;
      END
   END n_80905

   PIN n_80956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.69 61.277 48.718 61.44 ;
      END
   END n_80956

   PIN n_81032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.338 61.277 76.366 61.44 ;
      END
   END n_81032

   PIN n_81118
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.186 61.358 91.214 61.44 ;
      END
   END n_81118

   PIN n_81188
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.962 61.277 94.99 61.44 ;
      END
   END n_81188

   PIN n_81261
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.77 61.277 94.798 61.44 ;
      END
   END n_81261

   PIN n_81264
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.146 0.163 12.174 ;
      END
   END n_81264

   PIN n_81273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.066 0.0 14.094 0.163 ;
      END
   END n_81273

   PIN n_81298
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.09 61.277 23.118 61.44 ;
      END
   END n_81298

   PIN n_81301
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.442 61.277 99.47 61.44 ;
      END
   END n_81301

   PIN n_81360
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.586 61.277 17.614 61.44 ;
      END
   END n_81360

   PIN n_81395
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.122 61.277 91.15 61.44 ;
      END
   END n_81395

   PIN n_81420
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.41 0.082 7.438 ;
      END
   END n_81420

   PIN n_81431
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.09 0.163 7.118 ;
      END
   END n_81431

   PIN n_81462
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.674 0.163 18.702 ;
      END
   END n_81462

   PIN n_81477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.994 61.277 91.022 61.44 ;
      END
   END n_81477

   PIN n_81478
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.93 61.277 90.958 61.44 ;
      END
   END n_81478

   PIN n_81503
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.082 0.163 12.11 ;
      END
   END n_81503

   PIN n_81504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.538 0.163 7.566 ;
      END
   END n_81504

   PIN n_81590
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 73.266 61.277 73.294 61.44 ;
      END
   END n_81590

   PIN n_81626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.338 0.163 12.366 ;
      END
   END n_81626

   PIN n_81646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.682 61.277 109.71 61.44 ;
      END
   END n_81646

   PIN n_81668
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.162 0.163 2.19 ;
      END
   END n_81668

   PIN n_81761
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.986 0.163 8.014 ;
      END
   END n_81761

   PIN n_81776
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.018 61.277 76.046 61.44 ;
      END
   END n_81776

   PIN n_81799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.018 0.163 12.046 ;
      END
   END n_81799

   PIN n_81886
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.378 61.277 91.406 61.44 ;
      END
   END n_81886

   PIN n_81905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.97 61.277 97.998 61.44 ;
      END
   END n_81905

   PIN n_81907
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.578 61.277 94.606 61.44 ;
      END
   END n_81907

   PIN n_81908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.514 61.277 94.542 61.44 ;
      END
   END n_81908

   PIN n_81955
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.922 0.163 7.95 ;
      END
   END n_81955

   PIN n_82085
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.682 61.277 101.71 61.44 ;
      END
   END n_82085

   PIN n_82109
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.794 0.163 7.822 ;
      END
   END n_82109

   PIN n_82147
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.954 0.163 11.982 ;
      END
   END n_82147

   PIN n_82168
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.434 0.163 16.462 ;
      END
   END n_82168

   PIN n_82173
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.986 61.277 104.014 61.44 ;
      END
   END n_82173

   PIN n_82174
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.49 61.277 77.518 61.44 ;
      END
   END n_82174

   PIN n_82178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.738 61.277 90.766 61.44 ;
      END
   END n_82178

   PIN n_82215
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.37 0.163 16.398 ;
      END
   END n_82215

   PIN n_82244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.442 61.277 83.47 61.44 ;
      END
   END n_82244

   PIN n_82268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.442 61.277 91.47 61.44 ;
      END
   END n_82268

   PIN n_82282
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.058 0.163 11.086 ;
      END
   END n_82282

   PIN n_82287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.73 0.163 7.758 ;
      END
   END n_82287

   PIN n_82291
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.778 0.0 17.806 0.163 ;
      END
   END n_82291

   PIN n_82311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.09 61.277 95.118 61.44 ;
      END
   END n_82311

   PIN n_82329
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.89 0.163 11.918 ;
      END
   END n_82329

   PIN n_82352
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.474 61.277 79.502 61.44 ;
      END
   END n_82352

   PIN n_82357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.73 0.0 15.758 0.163 ;
      END
   END n_82357

   PIN n_82374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.05 0.163 8.078 ;
      END
   END n_82374

   PIN n_82375
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.618 61.277 21.646 61.44 ;
      END
   END n_82375

   PIN n_82412
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.65 61.277 105.678 61.44 ;
      END
   END n_82412

   PIN n_82417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.706 61.277 94.734 61.44 ;
      END
   END n_82417

   PIN n_82424
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.218 61.277 111.246 61.44 ;
      END
   END n_82424

   PIN n_82432
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.154 61.277 95.182 61.44 ;
      END
   END n_82432

   PIN n_82451
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.914 61.277 28.942 61.44 ;
      END
   END n_82451

   PIN n_82505
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.61 61.277 18.638 61.44 ;
      END
   END n_82505

   PIN n_82562
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.85 61.277 100.878 61.44 ;
      END
   END n_82562

   PIN n_82586
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.378 61.277 83.406 61.44 ;
      END
   END n_82586

   PIN n_82645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 26.866 0.163 26.894 ;
      END
   END n_82645

   PIN n_82650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.05 61.277 96.078 61.44 ;
      END
   END n_82650

   PIN n_82678
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.306 61.277 112.334 61.44 ;
      END
   END n_82678

   PIN n_82679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.138 61.277 25.166 61.44 ;
      END
   END n_82679

   PIN n_82698
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.45 0.163 30.478 ;
      END
   END n_82698

   PIN n_82738
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.17 61.277 29.198 61.44 ;
      END
   END n_82738

   PIN n_82745
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.098 61.277 26.126 61.44 ;
      END
   END n_82745

   PIN n_82764
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.162 61.277 26.19 61.44 ;
      END
   END n_82764

   PIN n_82769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.418 61.277 90.446 61.44 ;
      END
   END n_82769

   PIN n_82770
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.506 61.277 83.534 61.44 ;
      END
   END n_82770

   PIN n_83142
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.874 61.277 69.902 61.44 ;
      END
   END n_83142

   PIN n_83215
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 129.33 61.277 129.358 61.44 ;
      END
   END n_83215

   PIN n_84346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.402 61.277 132.43 61.44 ;
      END
   END n_84346

   PIN n_84639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.17 61.277 133.198 61.44 ;
      END
   END n_84639

   PIN n_84673
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.594 61.277 140.622 61.44 ;
      END
   END n_84673

   PIN n_84781
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 127.026 61.277 127.054 61.44 ;
      END
   END n_84781

   PIN n_84844
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.066 61.277 110.094 61.44 ;
      END
   END n_84844

   PIN n_99925
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.834 61.277 86.862 61.44 ;
      END
   END n_99925

   PIN stage2_out_3228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.738 61.277 2.766 61.44 ;
      END
   END stage2_out_3228

   PIN stage2_out_3231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.186 0.163 59.214 ;
      END
   END stage2_out_3231

   PIN stage2_out_3237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.522 0.163 49.55 ;
      END
   END stage2_out_3237

   PIN stage2_out_3238
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.354 61.277 10.382 61.44 ;
      END
   END stage2_out_3238

   PIN stage2_out_3262
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.714 61.277 25.742 61.44 ;
      END
   END stage2_out_3262

   PIN u1_L14_20_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.402 0.163 44.43 ;
      END
   END u1_L14_20_

   PIN u1_R13_16_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.922 0.163 39.95 ;
      END
   END u1_R13_16_

   PIN u1_R13_29_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.122 0.163 59.15 ;
      END
   END u1_R13_29_

   PIN u1_R13_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.002 0.163 54.03 ;
      END
   END u1_R13_6_

   PIN u2_IP_32_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.25 0.163 59.278 ;
      END
   END u2_IP_32_

   PIN u2_IP_64__1271
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.05 61.277 32.078 61.44 ;
      END
   END u2_IP_64__1271

   PIN u2_IP_64__1272
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.682 61.277 45.71 61.44 ;
      END
   END u2_IP_64__1272

   PIN u2_IP_64__1273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.162 61.277 34.19 61.44 ;
      END
   END u2_IP_64__1273

   PIN u2_IP_64__1278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.098 61.277 18.126 61.44 ;
      END
   END u2_IP_64__1278

   PIN u2_IP_64__1280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.49 61.277 37.518 61.44 ;
      END
   END u2_IP_64__1280

   PIN u2_IP_64__1282
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.25 61.277 3.278 61.44 ;
      END
   END u2_IP_64__1282

   PIN u2_IP_64__1286
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.81 61.277 21.838 61.44 ;
      END
   END u2_IP_64__1286

   PIN u2_L0_26_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.338 61.277 52.366 61.44 ;
      END
   END u2_L0_26_

   PIN u2_L0_31_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.21 61.277 60.238 61.44 ;
      END
   END u2_L0_31_

   PIN u2_L0_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.858 61.277 63.886 61.44 ;
      END
   END u2_L0_7_

   PIN u2_L0_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.026 61.277 79.054 61.44 ;
      END
   END u2_L0_9_

   PIN u2_L0_reg_10__Q
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.818 61.277 40.846 61.44 ;
      END
   END u2_L0_reg_10__Q

   PIN u2_L10_27_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.858 61.277 71.886 61.44 ;
      END
   END u2_L10_27_

   PIN u2_L10_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.866 61.277 82.894 61.44 ;
      END
   END u2_L10_5_

   PIN u2_L1_23_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.202 61.277 25.23 61.44 ;
      END
   END u2_L1_23_

   PIN u2_L1_28_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.922 61.277 71.95 61.44 ;
      END
   END u2_L1_28_

   PIN u2_L1_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.482 0.163 26.51 ;
      END
   END u2_L1_9_

   PIN u2_L1_reg_14__Q
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.874 61.277 29.902 61.44 ;
      END
   END u2_L1_reg_14__Q

   PIN u2_L2_18_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.786 61.277 44.814 61.44 ;
      END
   END u2_L2_18_

   PIN u2_R0_23_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.466 61.277 28.494 61.44 ;
      END
   END u2_R0_23_

   PIN u2_R0_25_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.21 61.277 36.238 61.44 ;
      END
   END u2_R0_25_

   PIN u2_R0_26_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.818 61.277 64.846 61.44 ;
      END
   END u2_R0_26_

   PIN u2_R0_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.37 61.277 152.398 61.44 ;
      END
   END u2_R0_5_

   PIN u2_R11_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.09 61.277 119.118 61.44 ;
      END
   END u2_R11_15_

   PIN u2_R11_21_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.05 61.277 112.078 61.44 ;
      END
   END u2_R11_21_

   PIN u2_R11_27_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.786 61.277 116.814 61.44 ;
      END
   END u2_R11_27_

   PIN u2_R12_22_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 156.274 61.277 156.302 61.44 ;
      END
   END u2_R12_22_

   PIN u2_R12_28_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.858 61.277 63.886 61.44 ;
      END
   END u2_R12_28_

   PIN u2_R13_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.53 61.277 52.558 61.44 ;
      END
   END u2_R13_5_

   PIN u2_R1_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.402 61.277 52.43 61.44 ;
      END
   END u2_R1_14_

   PIN u2_R1_30_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.194 61.277 54.222 61.44 ;
      END
   END u2_R1_30_

   PIN u2_R2_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.538 61.277 71.566 61.44 ;
      END
   END u2_R2_1_

   PIN u2_R2_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.682 61.277 21.71 61.44 ;
      END
   END u2_R2_3_

   PIN u2_R2_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.762 61.277 67.79 61.44 ;
      END
   END u2_R2_6_

   PIN u2_R2_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.514 61.277 118.542 61.44 ;
      END
   END u2_R2_7_

   PIN u2_key_r_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.018 61.277 60.046 61.44 ;
      END
   END u2_key_r_2_

   PIN u2_key_r_35_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.93 61.277 82.958 61.44 ;
      END
   END u2_key_r_35_

   PIN u2_key_r_55_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.562 61.277 56.59 61.44 ;
      END
   END u2_key_r_55_

   PIN u2_key_r_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.49 61.277 45.518 61.44 ;
      END
   END u2_key_r_5_

   PIN u2_uk_K_r_241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.922 61.277 71.95 61.44 ;
      END
   END u2_uk_K_r_241

   PIN u2_uk_K_r_270
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 61.277 25.614 61.44 ;
      END
   END u2_uk_K_r_270

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 167.36 61.44 ;
      LAYER V1 ;
         RECT 0.0 0.0 167.36 61.44 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 167.36 61.44 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 167.36 61.44 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 167.36 61.44 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 167.36 61.44 ;
      LAYER M1 ;
         RECT 0.0 0.0 167.36 61.44 ;
   END
END h2_mgc_des_perf_a

MACRO h1_mgc_des_perf_a
   CLASS BLOCK ;
   FOREIGN h1 ;
   ORIGIN 0 0 ;
   SIZE 106.624 BY 60.16 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1117_n_85315
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.234 59.997 93.262 60.16 ;
      END
   END FE_OFN1117_n_85315

   PIN FE_OFN1131_n_83717
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.258 106.624 46.286 ;
      END
   END FE_OFN1131_n_83717

   PIN FE_OFN1447_n_87131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.546 59.997 98.574 60.16 ;
      END
   END FE_OFN1447_n_87131

   PIN FE_OFN171_n_88228
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.842 59.997 81.87 60.16 ;
      END
   END FE_OFN171_n_88228

   PIN FE_OFN177_n_87818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.706 59.997 86.734 60.16 ;
      END
   END FE_OFN177_n_87818

   PIN FE_OFN183_n_87238
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.122 59.997 75.15 60.16 ;
      END
   END FE_OFN183_n_87238

   PIN FE_OFN2079_n_83196
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.914 59.997 100.942 60.16 ;
      END
   END FE_OFN2079_n_83196

   PIN FE_OFN2128_n_87090
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.97 59.997 81.998 60.16 ;
      END
   END FE_OFN2128_n_87090

   PIN FE_OFN2671_n_16014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 46.322 106.624 46.35 ;
      END
   END FE_OFN2671_n_16014

   PIN FE_OFN2969_n_15130
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.85 59.997 100.878 60.16 ;
      END
   END FE_OFN2969_n_15130

   PIN FE_OFN4075_n_84990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.45 59.997 102.478 60.16 ;
      END
   END FE_OFN4075_n_84990

   PIN g209359_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.962 59.997 62.99 60.16 ;
      END
   END g209359_p

   PIN g210571_p1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.906 59.997 81.934 60.16 ;
      END
   END g210571_p1

   PIN g210641_p2
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.554 59.997 93.582 60.16 ;
      END
   END g210641_p2

   PIN g210835_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.258 59.997 86.286 60.16 ;
      END
   END g210835_sb

   PIN g210889_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 30.322 106.624 30.35 ;
      END
   END g210889_p

   PIN g211048_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 31.026 106.624 31.054 ;
      END
   END g211048_p

   PIN g211616_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.418 106.624 50.446 ;
      END
   END g211616_p

   PIN g211975_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.97 59.997 81.998 60.16 ;
      END
   END g211975_db

   PIN g212677_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.41 59.997 95.438 60.16 ;
      END
   END g212677_p

   PIN g213393_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.906 59.997 97.934 60.16 ;
      END
   END g213393_p

   PIN g213779_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.258 59.997 102.286 60.16 ;
      END
   END g213779_p

   PIN g214217_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.746 59.997 101.774 60.16 ;
      END
   END g214217_db

   PIN g214217_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.834 59.997 102.862 60.16 ;
      END
   END g214217_sb

   PIN g214307_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.09 106.624 47.118 ;
      END
   END g214307_p

   PIN g214357_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.906 59.997 89.934 60.16 ;
      END
   END g214357_da

   PIN g215900_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.754 106.624 40.782 ;
      END
   END g215900_p

   PIN g305635_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.522 59.997 17.55 60.16 ;
      END
   END g305635_da

   PIN g305680_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.146 59.997 36.174 60.16 ;
      END
   END g305680_da

   PIN g305680_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.21 59.997 36.238 60.16 ;
      END
   END g305680_db

   PIN key_b_r_3__184
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.338 59.997 12.366 60.16 ;
      END
   END key_b_r_3__184

   PIN key_c_r_11__1306
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.218 59.997 31.246 60.16 ;
      END
   END key_c_r_11__1306

   PIN key_c_r_19__1727
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.314 59.997 59.342 60.16 ;
      END
   END key_c_r_19__1727

   PIN key_c_r_23__2371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.858 59.997 39.886 60.16 ;
      END
   END key_c_r_23__2371

   PIN key_c_r_28__2019
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.074 59.997 41.102 60.16 ;
      END
   END key_c_r_28__2019

   PIN key_c_r_29__2042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.578 0.0 102.606 0.163 ;
      END
   END key_c_r_29__2042

   PIN key_c_r_30__2096
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.026 59.997 55.054 60.16 ;
      END
   END key_c_r_30__2096

   PIN key_c_r_31__2167
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.53 59.997 92.558 60.16 ;
      END
   END key_c_r_31__2167

   PIN key_c_r_32__2208
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 3.762 106.624 3.79 ;
      END
   END key_c_r_32__2208

   PIN key_c_r_32__2234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.298 59.997 93.326 60.16 ;
      END
   END key_c_r_32__2234

   PIN key_c_r_33__17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.61 59.997 82.638 60.16 ;
      END
   END key_c_r_33__17_

   PIN key_c_r_33__29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 87.474 59.997 87.502 60.16 ;
      END
   END key_c_r_33__29_

   PIN key_c_r_33__41_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 54.002 106.624 54.03 ;
      END
   END key_c_r_33__41_

   PIN key_c_r_5__2758
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.018 59.997 12.046 60.16 ;
      END
   END key_c_r_5__2758

   PIN key_c_r_8__1129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.97 59.997 9.998 60.16 ;
      END
   END key_c_r_8__1129

   PIN n_117130
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.226 0.0 82.254 0.163 ;
      END
   END n_117130

   PIN n_117135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.066 0.0 86.094 0.163 ;
      END
   END n_117135

   PIN n_126115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 34.098 106.624 34.126 ;
      END
   END n_126115

   PIN n_15020
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.226 106.624 58.254 ;
      END
   END n_15020

   PIN n_15309
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.962 106.624 54.99 ;
      END
   END n_15309

   PIN n_15373
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.194 59.997 102.222 60.16 ;
      END
   END n_15373

   PIN n_15376
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.482 106.624 50.51 ;
      END
   END n_15376

   PIN n_15814
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.962 59.997 102.99 60.16 ;
      END
   END n_15814

   PIN n_16235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 46.386 106.624 46.414 ;
      END
   END n_16235

   PIN n_16236
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 55.026 106.624 55.054 ;
      END
   END n_16236

   PIN n_599
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.186 59.997 43.214 60.16 ;
      END
   END n_599

   PIN n_636
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.602 59.997 15.63 60.16 ;
      END
   END n_636

   PIN n_643
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.466 59.997 28.494 60.16 ;
      END
   END n_643

   PIN n_82873
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 35.89 106.624 35.918 ;
      END
   END n_82873

   PIN n_82885
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 42.162 106.624 42.19 ;
      END
   END n_82885

   PIN n_82988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.842 59.997 97.87 60.16 ;
      END
   END n_82988

   PIN n_83094
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.514 106.624 38.542 ;
      END
   END n_83094

   PIN n_83137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 47.09 106.624 47.118 ;
      END
   END n_83137

   PIN n_83203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.066 59.997 86.094 60.16 ;
      END
   END n_83203

   PIN n_83256
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 38.77 106.624 38.798 ;
      END
   END n_83256

   PIN n_83274
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.17 106.624 45.198 ;
      END
   END n_83274

   PIN n_83283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.218 106.624 39.246 ;
      END
   END n_83283

   PIN n_83296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.834 106.624 38.862 ;
      END
   END n_83296

   PIN n_83307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 11.506 106.624 11.534 ;
      END
   END n_83307

   PIN n_83371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 34.546 106.624 34.574 ;
      END
   END n_83371

   PIN n_83404
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 37.234 106.624 37.262 ;
      END
   END n_83404

   PIN n_83450
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.258 106.624 38.286 ;
      END
   END n_83450

   PIN n_83520
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.066 106.624 38.094 ;
      END
   END n_83520

   PIN n_83598
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.026 106.624 39.054 ;
      END
   END n_83598

   PIN n_83639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.97 106.624 49.998 ;
      END
   END n_83639

   PIN n_83663
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.642 106.624 38.67 ;
      END
   END n_83663

   PIN n_83674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 7.858 106.624 7.886 ;
      END
   END n_83674

   PIN n_83733
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 41.586 106.624 41.614 ;
      END
   END n_83733

   PIN n_83783
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.794 106.624 39.822 ;
      END
   END n_83783

   PIN n_83805
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.578 0.0 102.606 0.163 ;
      END
   END n_83805

   PIN n_83907
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.106 106.624 45.134 ;
      END
   END n_83907

   PIN n_83923
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 7.602 106.624 7.63 ;
      END
   END n_83923

   PIN n_83974
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.002 106.624 38.03 ;
      END
   END n_83974

   PIN n_84019
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.578 106.624 46.606 ;
      END
   END n_84019

   PIN n_84035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.578 106.624 38.606 ;
      END
   END n_84035

   PIN n_84063
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 41.65 106.624 41.678 ;
      END
   END n_84063

   PIN n_84124
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.898 106.624 38.926 ;
      END
   END n_84124

   PIN n_84128
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.114 106.624 40.142 ;
      END
   END n_84128

   PIN n_84129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.178 106.624 40.206 ;
      END
   END n_84129

   PIN n_84154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 34.418 106.624 34.446 ;
      END
   END n_84154

   PIN n_84252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.474 106.624 39.502 ;
      END
   END n_84252

   PIN n_84301
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 34.482 106.624 34.51 ;
      END
   END n_84301

   PIN n_84317
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 34.29 106.624 34.318 ;
      END
   END n_84317

   PIN n_84327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.962 106.624 38.99 ;
      END
   END n_84327

   PIN n_84402
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 38.834 106.624 38.862 ;
      END
   END n_84402

   PIN n_84435
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.978 106.624 45.006 ;
      END
   END n_84435

   PIN n_84440
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.818 106.624 40.846 ;
      END
   END n_84440

   PIN n_84544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 35.826 106.624 35.854 ;
      END
   END n_84544

   PIN n_84557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.858 106.624 39.886 ;
      END
   END n_84557

   PIN n_84593
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 42.482 106.624 42.51 ;
      END
   END n_84593

   PIN n_84597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 41.778 106.624 41.806 ;
      END
   END n_84597

   PIN n_84610
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 34.354 106.624 34.382 ;
      END
   END n_84610

   PIN n_84652
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.514 0.0 102.542 0.163 ;
      END
   END n_84652

   PIN n_84873
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.402 106.624 44.43 ;
      END
   END n_84873

   PIN n_84915
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.498 106.624 48.526 ;
      END
   END n_84915

   PIN n_84933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.362 106.624 45.39 ;
      END
   END n_84933

   PIN n_84971
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.466 106.624 44.494 ;
      END
   END n_84971

   PIN n_84986
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.034 106.624 50.062 ;
      END
   END n_84986

   PIN n_84988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.53 106.624 44.558 ;
      END
   END n_84988

   PIN n_84998
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.362 59.997 93.39 60.16 ;
      END
   END n_84998

   PIN n_84999
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.234 106.624 45.262 ;
      END
   END n_84999

   PIN n_85002
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 53.746 106.624 53.774 ;
      END
   END n_85002

   PIN n_85013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 47.602 106.624 47.63 ;
      END
   END n_85013

   PIN n_85031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.946 106.624 48.974 ;
      END
   END n_85031

   PIN n_85033
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.018 106.624 44.046 ;
      END
   END n_85033

   PIN n_85037
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.322 106.624 46.35 ;
      END
   END n_85037

   PIN n_85044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 37.298 106.624 37.326 ;
      END
   END n_85044

   PIN n_85059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.642 59.997 70.67 60.16 ;
      END
   END n_85059

   PIN n_85086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.578 59.997 102.606 60.16 ;
      END
   END n_85086

   PIN n_85103
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.194 59.997 94.222 60.16 ;
      END
   END n_85103

   PIN n_85147
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.778 59.997 97.806 60.16 ;
      END
   END n_85147

   PIN n_85176
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.226 59.997 90.254 60.16 ;
      END
   END n_85176

   PIN n_85187
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.386 106.624 46.414 ;
      END
   END n_85187

   PIN n_85208
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.562 106.624 48.59 ;
      END
   END n_85208

   PIN n_85249
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.426 59.997 93.454 60.16 ;
      END
   END n_85249

   PIN n_85270
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.162 59.997 98.19 60.16 ;
      END
   END n_85270

   PIN n_85275
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 50.098 106.624 50.126 ;
      END
   END n_85275

   PIN n_85344
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.542 49.65 106.624 49.678 ;
      END
   END n_85344

   PIN n_85378
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.61 59.997 82.638 60.16 ;
      END
   END n_85378

   PIN n_85405
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.778 59.997 89.806 60.16 ;
      END
   END n_85405

   PIN n_85406
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.258 59.997 94.286 60.16 ;
      END
   END n_85406

   PIN n_85475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.458 59.997 89.486 60.16 ;
      END
   END n_85475

   PIN n_85559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.45 106.624 54.478 ;
      END
   END n_85559

   PIN n_85684
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.45 60.078 86.478 60.16 ;
      END
   END n_85684

   PIN n_85696
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.29 59.997 90.318 60.16 ;
      END
   END n_85696

   PIN n_85699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.682 59.997 85.71 60.16 ;
      END
   END n_85699

   PIN n_85700
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.13 59.997 86.158 60.16 ;
      END
   END n_85700

   PIN n_85722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.842 106.624 49.87 ;
      END
   END n_85722

   PIN n_85818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.802 59.997 90.83 60.16 ;
      END
   END n_85818

   PIN n_85821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.97 59.997 89.998 60.16 ;
      END
   END n_85821

   PIN n_85842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.642 59.997 86.67 60.16 ;
      END
   END n_85842

   PIN n_85870
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.522 106.624 49.55 ;
      END
   END n_85870

   PIN n_85877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 53.874 106.624 53.902 ;
      END
   END n_85877

   PIN n_85878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 53.938 106.624 53.966 ;
      END
   END n_85878

   PIN n_85879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 53.682 106.624 53.71 ;
      END
   END n_85879

   PIN n_85946
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.986 59.997 72.014 60.16 ;
      END
   END n_85946

   PIN n_85967
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.458 106.624 49.486 ;
      END
   END n_85967

   PIN n_85970
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.49 59.997 93.518 60.16 ;
      END
   END n_85970

   PIN n_85991
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.97 106.624 49.998 ;
      END
   END n_85991

   PIN n_86002
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.29 106.624 58.318 ;
      END
   END n_86002

   PIN n_86110
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.898 59.997 86.926 60.16 ;
      END
   END n_86110

   PIN n_86119
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.066 59.997 86.094 60.16 ;
      END
   END n_86119

   PIN n_86129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.33 106.624 49.358 ;
      END
   END n_86129

   PIN n_86135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.674 59.997 90.702 60.16 ;
      END
   END n_86135

   PIN n_86142
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 57.97 106.624 57.998 ;
      END
   END n_86142

   PIN n_86146
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.354 106.624 58.382 ;
      END
   END n_86146

   PIN n_86151
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.362 106.624 45.39 ;
      END
   END n_86151

   PIN n_86152
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.554 59.997 93.582 60.16 ;
      END
   END n_86152

   PIN n_86238
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.13 59.997 86.158 60.16 ;
      END
   END n_86238

   PIN n_86246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.77 59.997 86.798 60.16 ;
      END
   END n_86246

   PIN n_86249
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.266 106.624 49.294 ;
      END
   END n_86249

   PIN n_86258
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.514 106.624 54.542 ;
      END
   END n_86258

   PIN n_86296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.002 106.624 54.03 ;
      END
   END n_86296

   PIN n_86305
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 55.09 106.624 55.118 ;
      END
   END n_86305

   PIN n_86355
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 35.122 106.624 35.15 ;
      END
   END n_86355

   PIN n_86362
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.618 59.997 93.646 60.16 ;
      END
   END n_86362

   PIN n_86364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.586 59.997 97.614 60.16 ;
      END
   END n_86364

   PIN n_86365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.482 60.078 82.51 60.16 ;
      END
   END n_86365

   PIN n_86383
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 53.938 106.624 53.966 ;
      END
   END n_86383

   PIN n_86431
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.418 106.624 58.446 ;
      END
   END n_86431

   PIN n_86433
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 33.202 106.624 33.23 ;
      END
   END n_86433

   PIN n_86440
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.034 59.997 90.062 60.16 ;
      END
   END n_86440

   PIN n_86479
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.49 59.997 93.518 60.16 ;
      END
   END n_86479

   PIN n_86494
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.522 59.997 89.55 60.16 ;
      END
   END n_86494

   PIN n_86540
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.258 59.997 94.286 60.16 ;
      END
   END n_86540

   PIN n_86551
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 55.154 106.624 55.182 ;
      END
   END n_86551

   PIN n_86592
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.194 59.997 86.222 60.16 ;
      END
   END n_86592

   PIN n_86600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.034 59.997 82.062 60.16 ;
      END
   END n_86600

   PIN n_86621
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.026 59.997 63.054 60.16 ;
      END
   END n_86621

   PIN n_86643
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.986 59.997 96.014 60.16 ;
      END
   END n_86643

   PIN n_86645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 53.746 106.624 53.774 ;
      END
   END n_86645

   PIN n_86646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.346 59.997 95.374 60.16 ;
      END
   END n_86646

   PIN n_86674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.09 59.997 63.118 60.16 ;
      END
   END n_86674

   PIN n_86688
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.65 59.997 97.678 60.16 ;
      END
   END n_86688

   PIN n_86724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.242 59.997 96.27 60.16 ;
      END
   END n_86724

   PIN n_86745
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.026 59.997 63.054 60.16 ;
      END
   END n_86745

   PIN n_86793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 42.546 106.624 42.574 ;
      END
   END n_86793

   PIN n_86805
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.874 59.997 93.902 60.16 ;
      END
   END n_86805

   PIN n_86808
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 34.226 106.624 34.254 ;
      END
   END n_86808

   PIN n_86828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 50.162 106.624 50.19 ;
      END
   END n_86828

   PIN n_86842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.01 106.624 49.038 ;
      END
   END n_86842

   PIN n_86858
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.746 106.624 45.774 ;
      END
   END n_86858

   PIN n_87007
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.098 106.624 50.126 ;
      END
   END n_87007

   PIN n_87056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.73 106.624 47.758 ;
      END
   END n_87056

   PIN n_87144
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.994 59.997 75.022 60.16 ;
      END
   END n_87144

   PIN n_87202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.642 59.997 94.67 60.16 ;
      END
   END n_87202

   PIN n_87212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.354 59.997 90.382 60.16 ;
      END
   END n_87212

   PIN n_87219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.542 22.898 106.624 22.926 ;
      END
   END n_87219

   PIN n_87221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.122 59.997 59.15 60.16 ;
      END
   END n_87221

   PIN n_87239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.642 59.997 78.67 60.16 ;
      END
   END n_87239

   PIN n_87240
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.034 59.997 82.062 60.16 ;
      END
   END n_87240

   PIN n_87294
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.546 59.997 74.574 60.16 ;
      END
   END n_87294

   PIN n_87311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.898 60.078 78.926 60.16 ;
      END
   END n_87311

   PIN n_87321
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 31.73 106.624 31.758 ;
      END
   END n_87321

   PIN n_87330
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.602 59.997 47.63 60.16 ;
      END
   END n_87330

   PIN n_87336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.834 59.997 86.862 60.16 ;
      END
   END n_87336

   PIN n_87368
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.738 59.997 82.766 60.16 ;
      END
   END n_87368

   PIN n_87394
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.386 59.997 94.414 60.16 ;
      END
   END n_87394

   PIN n_87399
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.61 59.997 74.638 60.16 ;
      END
   END n_87399

   PIN n_87412
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.058 59.997 75.086 60.16 ;
      END
   END n_87412

   PIN n_87421
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.578 59.997 78.606 60.16 ;
      END
   END n_87421

   PIN n_87424
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 22.066 106.624 22.094 ;
      END
   END n_87424

   PIN n_87472
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.542 47.346 106.624 47.374 ;
      END
   END n_87472

   PIN n_87486
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 22.13 106.624 22.158 ;
      END
   END n_87486

   PIN n_87498
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.77 59.997 78.798 60.16 ;
      END
   END n_87498

   PIN n_87530
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.058 59.997 75.086 60.16 ;
      END
   END n_87530

   PIN n_87556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.706 59.997 78.734 60.16 ;
      END
   END n_87556

   PIN n_87572
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.29 59.997 74.318 60.16 ;
      END
   END n_87572

   PIN n_87580
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.322 59.997 94.35 60.16 ;
      END
   END n_87580

   PIN n_87586
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 72.05 59.997 72.078 60.16 ;
      END
   END n_87586

   PIN n_87593
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 30.13 106.624 30.158 ;
      END
   END n_87593

   PIN n_87600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.098 59.997 82.126 60.16 ;
      END
   END n_87600

   PIN n_87616
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.194 59.997 86.222 60.16 ;
      END
   END n_87616

   PIN n_87642
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 22.194 106.624 22.222 ;
      END
   END n_87642

   PIN n_87644
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.226 59.997 82.254 60.16 ;
      END
   END n_87644

   PIN n_87648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.922 59.997 39.95 60.16 ;
      END
   END n_87648

   PIN n_87657
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 30.194 106.624 30.222 ;
      END
   END n_87657

   PIN n_87697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.514 60.078 94.542 60.16 ;
      END
   END n_87697

   PIN n_87745
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.378 59.997 91.406 60.16 ;
      END
   END n_87745

   PIN n_87752
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.098 59.997 90.126 60.16 ;
      END
   END n_87752

   PIN n_87753
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.322 59.997 86.35 60.16 ;
      END
   END n_87753

   PIN n_87757
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.226 59.997 98.254 60.16 ;
      END
   END n_87757

   PIN n_87789
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.282 59.997 55.31 60.16 ;
      END
   END n_87789

   PIN n_87794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.938 59.997 93.966 60.16 ;
      END
   END n_87794

   PIN n_87812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.674 59.997 74.702 60.16 ;
      END
   END n_87812

   PIN n_87816
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.034 59.997 98.062 60.16 ;
      END
   END n_87816

   PIN n_87818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 27.186 106.624 27.214 ;
      END
   END n_87818

   PIN n_87821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.77 59.997 70.798 60.16 ;
      END
   END n_87821

   PIN n_87839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.706 59.997 70.734 60.16 ;
      END
   END n_87839

   PIN n_87875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.674 59.997 82.702 60.16 ;
      END
   END n_87875

   PIN n_87932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.162 59.997 82.19 60.16 ;
      END
   END n_87932

   PIN n_87934
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.542 41.778 106.624 41.806 ;
      END
   END n_87934

   PIN n_87935
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.93 59.997 66.958 60.16 ;
      END
   END n_87935

   PIN n_87944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 72.114 59.997 72.142 60.16 ;
      END
   END n_87944

   PIN n_87945
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.154 59.997 63.182 60.16 ;
      END
   END n_87945

   PIN n_87951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.354 59.997 82.382 60.16 ;
      END
   END n_87951

   PIN n_88028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.746 59.997 85.774 60.16 ;
      END
   END n_88028

   PIN n_88056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.554 59.997 101.582 60.16 ;
      END
   END n_88056

   PIN n_88065
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.25 59.997 91.278 60.16 ;
      END
   END n_88065

   PIN n_88067
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.026 59.997 103.054 60.16 ;
      END
   END n_88067

   PIN n_88085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.258 59.997 86.286 60.16 ;
      END
   END n_88085

   PIN n_88092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.162 59.997 90.19 60.16 ;
      END
   END n_88092

   PIN n_88094
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.938 59.997 93.966 60.16 ;
      END
   END n_88094

   PIN n_88111
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.898 59.997 78.926 60.16 ;
      END
   END n_88111

   PIN n_88115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.29 59.997 98.318 60.16 ;
      END
   END n_88115

   PIN n_88121
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.346 59.997 55.374 60.16 ;
      END
   END n_88121

   PIN n_88124
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.002 59.997 94.03 60.16 ;
      END
   END n_88124

   PIN n_88191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.618 106.624 45.646 ;
      END
   END n_88191

   PIN n_88200
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.81 59.997 85.838 60.16 ;
      END
   END n_88200

   PIN n_88216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.386 59.997 94.414 60.16 ;
      END
   END n_88216

   PIN n_88257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 28.402 106.624 28.43 ;
      END
   END n_88257

   PIN n_88341
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.81 59.997 101.838 60.16 ;
      END
   END n_88341

   PIN n_88342
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 31.666 106.624 31.694 ;
      END
   END n_88342

   PIN n_88348
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.066 59.997 94.094 60.16 ;
      END
   END n_88348

   PIN n_88351
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.802 59.997 82.83 60.16 ;
      END
   END n_88351

   PIN n_88352
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.322 59.997 86.35 60.16 ;
      END
   END n_88352

   PIN n_88358
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.586 59.997 89.614 60.16 ;
      END
   END n_88358

   PIN n_88359
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 31.09 106.624 31.118 ;
      END
   END n_88359

   PIN n_88383
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.874 59.997 85.902 60.16 ;
      END
   END n_88383

   PIN n_88433
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.618 59.997 93.646 60.16 ;
      END
   END n_88433

   PIN n_88466
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.418 59.997 82.446 60.16 ;
      END
   END n_88466

   PIN n_88505
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.098 59.997 82.126 60.16 ;
      END
   END n_88505

   PIN n_88508
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.162 59.997 82.19 60.16 ;
      END
   END n_88508

   PIN n_88519
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.65 59.997 89.678 60.16 ;
      END
   END n_88519

   PIN n_88570
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.386 59.997 78.414 60.16 ;
      END
   END n_88570

   PIN n_88591
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.226 59.997 82.254 60.16 ;
      END
   END n_88591

   PIN n_88603
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 32.306 106.624 32.334 ;
      END
   END n_88603

   PIN n_88633
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.322 59.997 102.35 60.16 ;
      END
   END n_88633

   PIN n_88640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.354 59.997 74.382 60.16 ;
      END
   END n_88640

   PIN n_88657
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.322 59.997 94.35 60.16 ;
      END
   END n_88657

   PIN n_88669
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.29 59.997 82.318 60.16 ;
      END
   END n_88669

   PIN n_88670
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.13 59.997 102.158 60.16 ;
      END
   END n_88670

   PIN n_88681
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.682 59.997 93.71 60.16 ;
      END
   END n_88681

   PIN n_88726
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.25 106.624 43.278 ;
      END
   END n_88726

   PIN n_88770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.098 59.997 98.126 60.16 ;
      END
   END n_88770

   PIN n_88771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.786 59.997 100.814 60.16 ;
      END
   END n_88771

   PIN n_88781
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.738 59.997 74.766 60.16 ;
      END
   END n_88781

   PIN n_88782
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.418 59.997 74.446 60.16 ;
      END
   END n_88782

   PIN n_88793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 42.482 106.624 42.51 ;
      END
   END n_88793

   PIN n_88815
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 19.122 106.624 19.15 ;
      END
   END n_88815

   PIN n_88816
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.97 59.997 97.998 60.16 ;
      END
   END n_88816

   PIN n_88842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.61 59.997 98.638 60.16 ;
      END
   END n_88842

   PIN n_88874
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 22.77 106.624 22.798 ;
      END
   END n_88874

   PIN n_88877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.714 59.997 97.742 60.16 ;
      END
   END n_88877

   PIN n_88897
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.882 106.624 40.91 ;
      END
   END n_88897

   PIN n_89163
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.21 59.997 100.238 60.16 ;
      END
   END n_89163

   PIN n_89299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.002 59.997 94.03 60.16 ;
      END
   END n_89299

   PIN n_89430
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.546 106.624 50.574 ;
      END
   END n_89430

   PIN n_89487
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.522 59.997 97.55 60.16 ;
      END
   END n_89487

   PIN n_89527
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.834 59.997 70.862 60.16 ;
      END
   END n_89527

   PIN n_89607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.642 106.624 46.67 ;
      END
   END n_89607

   PIN n_89612
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.186 59.997 99.214 60.16 ;
      END
   END n_89612

   PIN n_89671
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.506 59.997 99.534 60.16 ;
      END
   END n_89671

   PIN n_89743
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.338 106.624 44.366 ;
      END
   END n_89743

   PIN n_89790
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.658 59.997 100.686 60.16 ;
      END
   END n_89790

   PIN n_89829
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.674 59.997 98.702 60.16 ;
      END
   END n_89829

   PIN n_89924
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.482 106.624 58.51 ;
      END
   END n_89924

   PIN n_89926
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 53.81 106.624 53.838 ;
      END
   END n_89926

   PIN n_89927
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.938 59.997 85.966 60.16 ;
      END
   END n_89927

   PIN n_89999
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.554 59.997 101.582 60.16 ;
      END
   END n_89999

   PIN n_90006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 46.194 106.624 46.222 ;
      END
   END n_90006

   PIN n_90059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.162 59.997 98.19 60.16 ;
      END
   END n_90059

   PIN n_90215
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.066 59.997 94.094 60.16 ;
      END
   END n_90215

   PIN n_90279
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.122 59.997 99.15 60.16 ;
      END
   END n_90279

   PIN n_90333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.994 59.997 99.022 60.16 ;
      END
   END n_90333

   PIN n_90412
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.994 59.997 99.022 60.16 ;
      END
   END n_90412

   PIN n_90417
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.618 59.997 101.646 60.16 ;
      END
   END n_90417

   PIN n_90560
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.994 59.997 67.022 60.16 ;
      END
   END n_90560

   PIN n_90687
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.978 59.997 101.006 60.16 ;
      END
   END n_90687

   PIN n_90693
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.546 106.624 58.574 ;
      END
   END n_90693

   PIN n_90818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.698 106.624 43.726 ;
      END
   END n_90818

   PIN n_90859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.594 106.624 44.622 ;
      END
   END n_90859

   PIN u1_key_r_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.57 59.997 75.598 60.16 ;
      END
   END u1_key_r_2_

   PIN u1_key_r_30_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.442 59.997 91.47 60.16 ;
      END
   END u1_key_r_30_

   PIN u1_key_r_55_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.986 59.997 80.014 60.16 ;
      END
   END u1_key_r_55_

   PIN u2_L2_17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.658 106.624 44.686 ;
      END
   END u2_L2_17_

   PIN u2_L3_18_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.898 59.997 70.926 60.16 ;
      END
   END u2_L3_18_

   PIN u2_L3_reg_14__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.066 59.997 102.094 60.16 ;
      END
   END u2_L3_reg_14__Q

   PIN u2_L4_18_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.514 106.624 46.542 ;
      END
   END u2_L4_18_

   PIN u2_L4_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.634 106.624 43.662 ;
      END
   END u2_L4_28_

   PIN u2_L4_32_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.738 59.997 74.766 60.16 ;
      END
   END u2_L4_32_

   PIN u2_L4_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.482 59.997 74.51 60.16 ;
      END
   END u2_L4_8_

   PIN u2_L5_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.722 106.624 44.75 ;
      END
   END u2_L5_14_

   PIN u2_L5_30_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.002 59.997 102.03 60.16 ;
      END
   END u2_L5_30_

   PIN u2_L5_reg_12__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.786 106.624 44.814 ;
      END
   END u2_L5_reg_12__Q

   PIN u2_R3_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.746 0.0 93.774 0.163 ;
      END
   END u2_R3_1_

   PIN u2_R3_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.194 59.997 102.222 60.16 ;
      END
   END u2_R3_2_

   PIN u2_R3_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.946 106.624 40.974 ;
      END
   END u2_R3_7_

   PIN u2_R4_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.354 59.997 82.382 60.16 ;
      END
   END u2_R4_13_

   PIN u2_R4_22_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.906 106.624 49.934 ;
      END
   END u2_R4_22_

   PIN u2_R4_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.61 106.624 58.638 ;
      END
   END u2_R4_23_

   PIN u2_R4_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.386 59.997 86.414 60.16 ;
      END
   END u2_R4_28_

   PIN u2_R4_29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.45 106.624 46.478 ;
      END
   END u2_R4_29_

   PIN u2_R4_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.746 59.997 93.774 60.16 ;
      END
   END u2_R4_3_

   PIN u2_R5_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.13 106.624 38.158 ;
      END
   END u2_R5_12_

   PIN u2_R5_29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 37.362 106.624 37.39 ;
      END
   END u2_R5_29_

   PIN u2_R5_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 19.186 106.624 19.214 ;
      END
   END u2_R5_4_

   PIN u2_key_r_21_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.026 59.997 71.054 60.16 ;
      END
   END u2_key_r_21_

   PIN u2_uk_K_r_530
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.274 106.624 44.302 ;
      END
   END u2_uk_K_r_530

   PIN FE_OFN1065_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.106 60.078 93.134 60.16 ;
      END
   END FE_OFN1065_n_116

   PIN FE_OFN1130_n_82876
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 42.546 106.624 42.574 ;
      END
   END FE_OFN1130_n_82876

   PIN FE_OFN1354_n_88664
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.33 106.624 49.358 ;
      END
   END FE_OFN1354_n_88664

   PIN FE_OFN1476_n_15154
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.522 106.624 41.55 ;
      END
   END FE_OFN1476_n_15154

   PIN FE_OFN1597_n_16688
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 37.042 106.624 37.07 ;
      END
   END FE_OFN1597_n_16688

   PIN FE_OFN176_n_87818
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 27.122 106.624 27.15 ;
      END
   END FE_OFN176_n_87818

   PIN FE_OFN1837_n_16002
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 41.842 106.624 41.87 ;
      END
   END FE_OFN1837_n_16002

   PIN FE_OFN1909_n_85016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.026 106.624 47.054 ;
      END
   END FE_OFN1909_n_85016

   PIN FE_OFN2000_n_84960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.138 106.624 41.166 ;
      END
   END FE_OFN2000_n_84960

   PIN FE_OFN2127_n_87090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.226 59.997 74.254 60.16 ;
      END
   END FE_OFN2127_n_87090

   PIN FE_OFN2410_n_82958
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 57.586 106.624 57.614 ;
      END
   END FE_OFN2410_n_82958

   PIN FE_OFN2514_n_82929
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.542 39.666 106.624 39.694 ;
      END
   END FE_OFN2514_n_82929

   PIN FE_OFN2809_n_16012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 57.906 106.624 57.934 ;
      END
   END FE_OFN2809_n_16012

   PIN FE_OFN2888_n_16011
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.53 59.997 100.558 60.16 ;
      END
   END FE_OFN2888_n_16011

   PIN FE_OFN3132_n_16013
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 43.122 106.624 43.15 ;
      END
   END FE_OFN3132_n_16013

   PIN FE_OFN3225_n_15131
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.962 106.624 46.99 ;
      END
   END FE_OFN3225_n_15131

   PIN FE_OFN3320_n_500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.986 60.078 16.014 60.16 ;
      END
   END FE_OFN3320_n_500

   PIN FE_OFN3436_n_89910
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.378 59.997 99.406 60.16 ;
      END
   END FE_OFN3436_n_89910

   PIN FE_OFN3698_n_16007
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.354 59.997 98.382 60.16 ;
      END
   END FE_OFN3698_n_16007

   PIN FE_OFN4024_n_85019
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 42.802 106.624 42.83 ;
      END
   END FE_OFN4024_n_85019

   PIN FE_OFN4400_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.542 49.586 106.624 49.614 ;
      END
   END FE_OFN4400_decrypt

   PIN FE_OFN4722_n_500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.61 60.078 74.638 60.16 ;
      END
   END FE_OFN4722_n_500

   PIN FE_OFN4816_n_16014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.898 106.624 54.926 ;
      END
   END FE_OFN4816_n_16014

   PIN FE_OFN872_n_84986
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.162 106.624 50.19 ;
      END
   END FE_OFN872_n_84986

   PIN g210626_p1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.354 59.997 74.382 60.16 ;
      END
   END g210626_p1

   PIN g210918_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.874 59.997 101.902 60.16 ;
      END
   END g210918_p

   PIN g211000_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.866 59.997 66.894 60.16 ;
      END
   END g211000_p

   PIN g211245_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.666 106.624 47.694 ;
      END
   END g211245_p

   PIN g211261_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 23.922 106.624 23.95 ;
      END
   END g211261_p

   PIN g211472_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.906 59.997 81.934 60.16 ;
      END
   END g211472_p

   PIN g211617_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.578 59.997 70.606 60.16 ;
      END
   END g211617_p

   PIN g211748_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.426 59.997 93.454 60.16 ;
      END
   END g211748_p

   PIN g212987_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.002 59.997 86.03 60.16 ;
      END
   END g212987_p

   PIN g214406_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.866 59.997 98.894 60.16 ;
      END
   END g214406_db

   PIN g214423_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.954 106.624 43.982 ;
      END
   END g214423_db

   PIN g214423_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.186 106.624 43.214 ;
      END
   END g214423_sb

   PIN g216122_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.194 106.624 46.222 ;
      END
   END g216122_sb

   PIN g216695_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.786 59.997 100.814 60.16 ;
      END
   END g216695_sb

   PIN g286480_p
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.834 106.624 54.862 ;
      END
   END g286480_p

   PIN g305627_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.65 59.997 17.678 60.16 ;
      END
   END g305627_sb

   PIN g305634_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.786 59.997 20.814 60.16 ;
      END
   END g305634_da

   PIN g305634_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.626 59.997 16.654 60.16 ;
      END
   END g305634_db

   PIN g305715_da
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.666 59.997 15.694 60.16 ;
      END
   END g305715_da

   PIN g321810_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.778 59.997 81.806 60.16 ;
      END
   END g321810_db

   PIN g321810_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.714 59.997 81.742 60.16 ;
      END
   END g321810_sb

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.542 42.29 106.624 42.318 ;
      END
   END ispd_clk

   PIN key1_17_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.586 59.997 17.614 60.16 ;
      END
   END key1_17_

   PIN key1_37_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.378 59.997 43.406 60.16 ;
      END
   END key1_37_

   PIN key1_39_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.482 59.997 74.51 60.16 ;
      END
   END key1_39_

   PIN key2_19_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.226 0.163 42.254 ;
      END
   END key2_19_

   PIN key3_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.45 59.997 14.478 60.16 ;
      END
   END key3_11_

   PIN key3_37_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.754 59.997 16.782 60.16 ;
      END
   END key3_37_

   PIN key3_39_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.418 59.997 74.446 60.16 ;
      END
   END key3_39_

   PIN key_b_r_15__880
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.026 59.997 47.054 60.16 ;
      END
   END key_b_r_15__880

   PIN key_b_r_16__2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.458 59.997 9.486 60.16 ;
      END
   END key_b_r_16__2_

   PIN key_b_r_16__30_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.042 59.997 13.07 60.16 ;
      END
   END key_b_r_16__30_

   PIN key_c_r_20__1782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.898 59.997 62.926 60.16 ;
      END
   END key_c_r_20__1782

   PIN key_c_r_21__1822
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.394 59.997 9.422 60.16 ;
      END
   END key_c_r_21__1822

   PIN key_c_r_27__1931
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.354 59.997 50.382 60.16 ;
      END
   END key_c_r_27__1931

   PIN key_c_r_27__1964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.082 59.997 36.11 60.16 ;
      END
   END key_c_r_27__1964

   PIN key_c_r_27__1966
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.018 59.997 36.046 60.16 ;
      END
   END key_c_r_27__1966

   PIN key_c_r_2__2648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.09 59.997 7.118 60.16 ;
      END
   END key_c_r_2__2648

   PIN key_c_r_30__2098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.69 59.997 24.718 60.16 ;
      END
   END key_c_r_30__2098

   PIN key_c_r_31__2162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.426 59.997 5.454 60.16 ;
      END
   END key_c_r_31__2162

   PIN key_c_r_31__2179
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.626 59.997 24.654 60.16 ;
      END
   END key_c_r_31__2179

   PIN key_c_r_32__2221
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.33 59.997 9.358 60.16 ;
      END
   END key_c_r_32__2221

   PIN key_c_r_32__2229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.562 59.997 24.59 60.16 ;
      END
   END key_c_r_32__2229

   PIN key_c_r_5__2791
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.266 59.997 9.294 60.16 ;
      END
   END key_c_r_5__2791

   PIN key_c_r_6__1019
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.426 59.997 5.454 60.16 ;
      END
   END key_c_r_6__1019

   PIN key_c_r_7__1051
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.714 59.997 33.742 60.16 ;
      END
   END key_c_r_7__1051

   PIN key_c_r_9__1177
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.274 59.997 36.302 60.16 ;
      END
   END key_c_r_9__1177

   PIN n_108924
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.938 59.997 85.966 60.16 ;
      END
   END n_108924

   PIN n_108925
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.65 59.997 81.678 60.16 ;
      END
   END n_108925

   PIN n_118831
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.714 59.997 97.742 60.16 ;
      END
   END n_118831

   PIN n_118867
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.866 59.997 66.894 60.16 ;
      END
   END n_118867

   PIN n_14583
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.162 106.624 58.19 ;
      END
   END n_14583

   PIN n_15021
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.89 106.624 43.918 ;
      END
   END n_15021

   PIN n_15130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.13 106.624 46.158 ;
      END
   END n_15130

   PIN n_15136
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.17 59.997 101.198 60.16 ;
      END
   END n_15136

   PIN n_15152
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.042 59.997 101.07 60.16 ;
      END
   END n_15152

   PIN n_15372
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.234 59.997 101.262 60.16 ;
      END
   END n_15372

   PIN n_15780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.77 106.624 54.798 ;
      END
   END n_15780

   PIN n_15789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.098 106.624 58.126 ;
      END
   END n_15789

   PIN n_15811
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.426 59.997 101.454 60.16 ;
      END
   END n_15811

   PIN n_15813
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.386 106.624 54.414 ;
      END
   END n_15813

   PIN n_15820
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.322 106.624 54.35 ;
      END
   END n_15820

   PIN n_15823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 57.842 106.624 57.87 ;
      END
   END n_15823

   PIN n_15989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.202 106.624 41.23 ;
      END
   END n_15989

   PIN n_16001
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.594 59.997 100.622 60.16 ;
      END
   END n_16001

   PIN n_16005
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 53.874 106.624 53.902 ;
      END
   END n_16005

   PIN n_16006
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.85 106.624 44.878 ;
      END
   END n_16006

   PIN n_16008
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.938 59.997 101.966 60.16 ;
      END
   END n_16008

   PIN n_16010
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 57.778 106.624 57.806 ;
      END
   END n_16010

   PIN n_16015
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.362 59.997 93.39 60.16 ;
      END
   END n_16015

   PIN n_16017
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.378 106.624 43.406 ;
      END
   END n_16017

   PIN n_16021
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.258 106.624 54.286 ;
      END
   END n_16021

   PIN n_16022
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 44.914 106.624 44.942 ;
      END
   END n_16022

   PIN n_16140
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 57.714 106.624 57.742 ;
      END
   END n_16140

   PIN n_16141
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.618 59.997 101.646 60.16 ;
      END
   END n_16141

   PIN n_16195
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.602 106.624 47.63 ;
      END
   END n_16195

   PIN n_16229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.81 106.624 45.838 ;
      END
   END n_16229

   PIN n_16233
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.386 59.997 102.414 60.16 ;
      END
   END n_16233

   PIN n_16511
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.802 59.997 98.83 60.16 ;
      END
   END n_16511

   PIN n_16677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 57.65 106.624 57.678 ;
      END
   END n_16677

   PIN n_16679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.218 106.624 47.246 ;
      END
   END n_16679

   PIN n_16680
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.322 59.997 102.35 60.16 ;
      END
   END n_16680

   PIN n_16684
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.482 59.997 98.51 60.16 ;
      END
   END n_16684

   PIN n_212558
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.842 59.997 81.87 60.16 ;
      END
   END n_212558

   PIN n_82772
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 42.034 106.624 42.062 ;
      END
   END n_82772

   PIN n_82780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.314 106.624 43.342 ;
      END
   END n_82780

   PIN n_82909
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.898 106.624 46.926 ;
      END
   END n_82909

   PIN n_83007
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.586 106.624 41.614 ;
      END
   END n_83007

   PIN n_83063
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 11.442 106.624 11.47 ;
      END
   END n_83063

   PIN n_83143
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 40.626 106.624 40.654 ;
      END
   END n_83143

   PIN n_83196
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 47.026 106.624 47.054 ;
      END
   END n_83196

   PIN n_83220
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.434 106.624 48.462 ;
      END
   END n_83220

   PIN n_83253
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.542 49.202 106.624 49.23 ;
      END
   END n_83253

   PIN n_83284
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.538 106.624 47.566 ;
      END
   END n_83284

   PIN n_83297
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 30.258 106.624 30.286 ;
      END
   END n_83297

   PIN n_83370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.09 106.624 39.118 ;
      END
   END n_83370

   PIN n_83394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.066 106.624 46.094 ;
      END
   END n_83394

   PIN n_83464
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.77 106.624 38.798 ;
      END
   END n_83464

   PIN n_83518
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 38.898 106.624 38.926 ;
      END
   END n_83518

   PIN n_83537
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.37 106.624 48.398 ;
      END
   END n_83537

   PIN n_83544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.49 106.624 45.518 ;
      END
   END n_83544

   PIN n_83637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.058 106.624 43.086 ;
      END
   END n_83637

   PIN n_83660
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.882 106.624 48.91 ;
      END
   END n_83660

   PIN n_83662
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 38.002 106.624 38.03 ;
      END
   END n_83662

   PIN n_83713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 41.714 106.624 41.742 ;
      END
   END n_83713

   PIN n_83717
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.002 106.624 46.03 ;
      END
   END n_83717

   PIN n_83770
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.154 106.624 39.182 ;
      END
   END n_83770

   PIN n_83804
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 3.826 106.624 3.854 ;
      END
   END n_83804

   PIN n_83818
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.298 106.624 45.326 ;
      END
   END n_83818

   PIN n_83848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.298 106.624 45.326 ;
      END
   END n_83848

   PIN n_83939
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.542 7.73 106.624 7.758 ;
      END
   END n_83939

   PIN n_83944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.346 106.624 39.374 ;
      END
   END n_83944

   PIN n_84141
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.834 106.624 46.862 ;
      END
   END n_84141

   PIN n_84142
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.586 0.0 97.614 0.163 ;
      END
   END n_84142

   PIN n_84180
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.69 106.624 40.718 ;
      END
   END n_84180

   PIN n_84307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.842 59.997 89.87 60.16 ;
      END
   END n_84307

   PIN n_84316
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 38.706 106.624 38.734 ;
      END
   END n_84316

   PIN n_84391
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.41 106.624 39.438 ;
      END
   END n_84391

   PIN n_84580
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.562 106.624 40.59 ;
      END
   END n_84580

   PIN n_84632
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.474 106.624 47.502 ;
      END
   END n_84632

   PIN n_84645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.05 106.624 40.078 ;
      END
   END n_84645

   PIN n_84646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.986 106.624 40.014 ;
      END
   END n_84646

   PIN n_84687
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.074 106.624 41.102 ;
      END
   END n_84687

   PIN n_84688
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.01 106.624 41.038 ;
      END
   END n_84688

   PIN n_84801
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.826 106.624 43.854 ;
      END
   END n_84801

   PIN n_84811
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 46.962 106.624 46.99 ;
      END
   END n_84811

   PIN n_84823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 40.562 106.624 40.59 ;
      END
   END n_84823

   PIN n_84840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 50.034 106.624 50.062 ;
      END
   END n_84840

   PIN n_84875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.282 106.624 39.31 ;
      END
   END n_84875

   PIN n_84895
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.898 59.997 102.926 60.16 ;
      END
   END n_84895

   PIN n_84903
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.506 106.624 43.534 ;
      END
   END n_84903

   PIN n_84918
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.682 59.997 101.71 60.16 ;
      END
   END n_84918

   PIN n_84940
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.77 106.624 46.798 ;
      END
   END n_84940

   PIN n_84990
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.45 59.997 102.478 60.16 ;
      END
   END n_84990

   PIN n_85014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.682 106.624 45.71 ;
      END
   END n_85014

   PIN n_85057
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.466 59.997 28.494 60.16 ;
      END
   END n_85057

   PIN n_85084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.554 106.624 45.582 ;
      END
   END n_85084

   PIN n_85194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 53.81 106.624 53.838 ;
      END
   END n_85194

   PIN n_85234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.874 59.997 85.902 60.16 ;
      END
   END n_85234

   PIN n_85248
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.738 59.997 90.766 60.16 ;
      END
   END n_85248

   PIN n_85335
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.034 59.997 98.062 60.16 ;
      END
   END n_85335

   PIN n_85437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.542 47.218 106.624 47.246 ;
      END
   END n_85437

   PIN n_85457
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.778 59.997 89.806 60.16 ;
      END
   END n_85457

   PIN n_85462
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.874 59.997 93.902 60.16 ;
      END
   END n_85462

   PIN n_85470
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.578 59.997 102.606 60.16 ;
      END
   END n_85470

   PIN n_85495
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.426 59.997 101.454 60.16 ;
      END
   END n_85495

   PIN n_85591
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.29 59.997 74.318 60.16 ;
      END
   END n_85591

   PIN n_85698
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 36.722 106.624 36.75 ;
      END
   END n_85698

   PIN n_85825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.714 59.997 89.742 60.16 ;
      END
   END n_85825

   PIN n_85840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.81 59.997 85.838 60.16 ;
      END
   END n_85840

   PIN n_85969
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.65 59.997 89.678 60.16 ;
      END
   END n_85969

   PIN n_85975
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.746 59.997 85.774 60.16 ;
      END
   END n_85975

   PIN n_86111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.682 59.997 85.71 60.16 ;
      END
   END n_86111

   PIN n_86144
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.906 106.624 49.934 ;
      END
   END n_86144

   PIN n_86164
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.706 106.624 54.734 ;
      END
   END n_86164

   PIN n_86241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.586 59.997 89.614 60.16 ;
      END
   END n_86241

   PIN n_86242
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.322 59.997 78.35 60.16 ;
      END
   END n_86242

   PIN n_86243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.81 59.997 93.838 60.16 ;
      END
   END n_86243

   PIN n_86295
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.194 106.624 54.222 ;
      END
   END n_86295

   PIN n_86457
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.13 106.624 54.158 ;
      END
   END n_86457

   PIN n_86466
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.778 106.624 49.806 ;
      END
   END n_86466

   PIN n_86468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 57.522 106.624 57.55 ;
      END
   END n_86468

   PIN n_86472
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.978 59.997 93.006 60.16 ;
      END
   END n_86472

   PIN n_86473
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.914 59.997 92.942 60.16 ;
      END
   END n_86473

   PIN n_86493
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.578 59.997 86.606 60.16 ;
      END
   END n_86493

   PIN n_86500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.618 59.997 85.646 60.16 ;
      END
   END n_86500

   PIN n_86542
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.066 106.624 54.094 ;
      END
   END n_86542

   PIN n_86577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.642 106.624 54.67 ;
      END
   END n_86577

   PIN n_86583
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.45 59.997 94.478 60.16 ;
      END
   END n_86583

   PIN n_86594
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.778 59.997 97.806 60.16 ;
      END
   END n_86594

   PIN n_86596
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.522 59.997 89.55 60.16 ;
      END
   END n_86596

   PIN n_86598
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.714 59.997 89.742 60.16 ;
      END
   END n_86598

   PIN n_86602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.818 106.624 48.846 ;
      END
   END n_86602

   PIN n_86605
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.554 59.997 85.582 60.16 ;
      END
   END n_86605

   PIN n_86618
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 54.578 106.624 54.606 ;
      END
   END n_86618

   PIN n_86641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.618 59.997 85.646 60.16 ;
      END
   END n_86641

   PIN n_86642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 49.394 106.624 49.422 ;
      END
   END n_86642

   PIN n_86644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.554 59.997 85.582 60.16 ;
      END
   END n_86644

   PIN n_86648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.106 106.624 45.134 ;
      END
   END n_86648

   PIN n_86690
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.33 59.997 97.358 60.16 ;
      END
   END n_86690

   PIN n_86691
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.298 59.997 93.326 60.16 ;
      END
   END n_86691

   PIN n_86696
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 42.802 106.624 42.83 ;
      END
   END n_86696

   PIN n_86750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.85 59.997 92.878 60.16 ;
      END
   END n_86750

   PIN n_86804
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.458 59.997 89.486 60.16 ;
      END
   END n_86804

   PIN n_86806
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.49 59.997 85.518 60.16 ;
      END
   END n_86806

   PIN n_86807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.234 59.997 93.262 60.16 ;
      END
   END n_86807

   PIN n_86815
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.642 59.997 102.67 60.16 ;
      END
   END n_86815

   PIN n_86816
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.706 59.997 102.734 60.16 ;
      END
   END n_86816

   PIN n_86829
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.394 59.997 89.422 60.16 ;
      END
   END n_86829

   PIN n_86839
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.434 59.997 96.462 60.16 ;
      END
   END n_86839

   PIN n_86843
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.938 106.624 45.966 ;
      END
   END n_86843

   PIN n_86851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 58.034 106.624 58.062 ;
      END
   END n_86851

   PIN n_86861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 37.17 106.624 37.198 ;
      END
   END n_86861

   PIN n_86969
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.994 59.997 75.022 60.16 ;
      END
   END n_86969

   PIN n_87008
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.122 106.624 43.15 ;
      END
   END n_87008

   PIN n_87034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.866 59.997 74.894 60.16 ;
      END
   END n_87034

   PIN n_87060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 27.442 106.624 27.47 ;
      END
   END n_87060

   PIN n_87145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 32.882 106.624 32.91 ;
      END
   END n_87145

   PIN n_87155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 29.042 106.624 29.07 ;
      END
   END n_87155

   PIN n_87159
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 30.962 106.624 30.99 ;
      END
   END n_87159

   PIN n_87178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.81 59.997 93.838 60.16 ;
      END
   END n_87178

   PIN n_87180
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.578 59.997 78.606 60.16 ;
      END
   END n_87180

   PIN n_87185
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.394 106.624 49.422 ;
      END
   END n_87185

   PIN n_87213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.97 106.624 41.998 ;
      END
   END n_87213

   PIN n_87230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.314 59.997 91.342 60.16 ;
      END
   END n_87230

   PIN n_87235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.354 106.624 50.382 ;
      END
   END n_87235

   PIN n_87275
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.154 106.624 47.182 ;
      END
   END n_87275

   PIN n_87293
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.546 59.997 82.574 60.16 ;
      END
   END n_87293

   PIN n_87322
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.258 59.997 78.286 60.16 ;
      END
   END n_87322

   PIN n_87328
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 31.282 106.624 31.31 ;
      END
   END n_87328

   PIN n_87329
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 30.514 106.624 30.542 ;
      END
   END n_87329

   PIN n_87354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.65 59.997 97.678 60.16 ;
      END
   END n_87354

   PIN n_87367
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.962 59.997 70.99 60.16 ;
      END
   END n_87367

   PIN n_87409
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.194 59.997 78.222 60.16 ;
      END
   END n_87409

   PIN n_87410
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.13 59.997 78.158 60.16 ;
      END
   END n_87410

   PIN n_87427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.906 59.997 97.934 60.16 ;
      END
   END n_87427

   PIN n_87453
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.194 59.997 94.222 60.16 ;
      END
   END n_87453

   PIN n_87468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.834 59.997 78.862 60.16 ;
      END
   END n_87468

   PIN n_87487
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.866 60.078 74.894 60.16 ;
      END
   END n_87487

   PIN n_87488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.426 59.997 85.454 60.16 ;
      END
   END n_87488

   PIN n_87493
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 29.682 106.624 29.71 ;
      END
   END n_87493

   PIN n_87500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.026 59.997 79.054 60.16 ;
      END
   END n_87500

   PIN n_87508
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.514 59.997 78.542 60.16 ;
      END
   END n_87508

   PIN n_87509
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.066 59.997 78.094 60.16 ;
      END
   END n_87509

   PIN n_87518
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.002 59.997 86.03 60.16 ;
      END
   END n_87518

   PIN n_87532
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.77 59.997 78.798 60.16 ;
      END
   END n_87532

   PIN n_87574
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.578 59.997 70.606 60.16 ;
      END
   END n_87574

   PIN n_87595
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.306 106.624 48.334 ;
      END
   END n_87595

   PIN n_87624
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.362 59.997 85.39 60.16 ;
      END
   END n_87624

   PIN n_87630
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.226 59.997 74.254 60.16 ;
      END
   END n_87630

   PIN n_87656
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.706 59.997 78.734 60.16 ;
      END
   END n_87656

   PIN n_87658
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.13 59.997 94.158 60.16 ;
      END
   END n_87658

   PIN n_87663
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.482 59.997 82.51 60.16 ;
      END
   END n_87663

   PIN n_87665
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.586 59.997 97.614 60.16 ;
      END
   END n_87665

   PIN n_87666
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.586 59.997 81.614 60.16 ;
      END
   END n_87666

   PIN n_87668
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 31.602 106.624 31.63 ;
      END
   END n_87668

   PIN n_87689
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.41 106.624 47.438 ;
      END
   END n_87689

   PIN n_87742
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.802 59.997 74.83 60.16 ;
      END
   END n_87742

   PIN n_87751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.514 59.997 78.542 60.16 ;
      END
   END n_87751

   PIN n_87756
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.842 59.997 97.87 60.16 ;
      END
   END n_87756

   PIN n_87776
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.754 106.624 48.782 ;
      END
   END n_87776

   PIN n_87779
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.45 59.997 78.478 60.16 ;
      END
   END n_87779

   PIN n_87782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.002 59.997 78.03 60.16 ;
      END
   END n_87782

   PIN n_87803
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 31.154 106.624 31.182 ;
      END
   END n_87803

   PIN n_87807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.802 59.997 66.83 60.16 ;
      END
   END n_87807

   PIN n_87810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.514 59.997 70.542 60.16 ;
      END
   END n_87810

   PIN n_87819
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.162 59.997 74.19 60.16 ;
      END
   END n_87819

   PIN n_87842
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.69 106.624 48.718 ;
      END
   END n_87842

   PIN n_87860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.45 59.997 70.478 60.16 ;
      END
   END n_87860

   PIN n_87863
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.29 59.997 82.318 60.16 ;
      END
   END n_87863

   PIN n_87872
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.298 59.997 85.326 60.16 ;
      END
   END n_87872

   PIN n_87884
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.162 59.997 74.19 60.16 ;
      END
   END n_87884

   PIN n_87897
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.834 59.997 62.862 60.16 ;
      END
   END n_87897

   PIN n_87911
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.57 106.624 43.598 ;
      END
   END n_87911

   PIN n_87937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.986 59.997 40.014 60.16 ;
      END
   END n_87937

   PIN n_87953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.29 106.624 50.318 ;
      END
   END n_87953

   PIN n_87954
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.874 106.624 45.902 ;
      END
   END n_87954

   PIN n_87964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.97 59.997 97.998 60.16 ;
      END
   END n_87964

   PIN n_87971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 22.002 106.624 22.03 ;
      END
   END n_87971

   PIN n_87976
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 32.242 106.624 32.27 ;
      END
   END n_87976

   PIN n_87986
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.394 59.997 89.422 60.16 ;
      END
   END n_87986

   PIN n_88058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.746 59.997 93.774 60.16 ;
      END
   END n_88058

   PIN n_88113
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.098 59.997 74.126 60.16 ;
      END
   END n_88113

   PIN n_88117
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 26.738 106.624 26.766 ;
      END
   END n_88117

   PIN n_88193
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.21 106.624 44.238 ;
      END
   END n_88193

   PIN n_88207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.45 59.997 78.478 60.16 ;
      END
   END n_88207

   PIN n_88213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.458 106.624 49.486 ;
      END
   END n_88213

   PIN n_88245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.234 59.997 85.262 60.16 ;
      END
   END n_88245

   PIN n_88254
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.234 106.624 45.262 ;
      END
   END n_88254

   PIN n_88256
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.002 59.997 102.03 60.16 ;
      END
   END n_88256

   PIN n_88259
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.066 59.997 102.094 60.16 ;
      END
   END n_88259

   PIN n_88261
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.17 59.997 93.198 60.16 ;
      END
   END n_88261

   PIN n_88265
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 44.082 106.624 44.11 ;
      END
   END n_88265

   PIN n_88318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.242 106.624 48.27 ;
      END
   END n_88318

   PIN n_88320
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.458 106.624 41.486 ;
      END
   END n_88320

   PIN n_88346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.81 106.624 45.838 ;
      END
   END n_88346

   PIN n_88381
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.386 59.997 70.414 60.16 ;
      END
   END n_88381

   PIN n_88397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.746 106.624 45.774 ;
      END
   END n_88397

   PIN n_88416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.106 59.997 93.134 60.16 ;
      END
   END n_88416

   PIN n_88417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.042 59.997 93.07 60.16 ;
      END
   END n_88417

   PIN n_88426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 48.626 106.624 48.654 ;
      END
   END n_88426

   PIN n_88428
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.842 106.624 49.87 ;
      END
   END n_88428

   PIN n_88454
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.074 106.624 49.102 ;
      END
   END n_88454

   PIN n_88468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.282 59.997 55.31 60.16 ;
      END
   END n_88468

   PIN n_88469
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.978 59.997 93.006 60.16 ;
      END
   END n_88469

   PIN n_88523
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.93 59.997 74.958 60.16 ;
      END
   END n_88523

   PIN n_88555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.17 106.624 45.198 ;
      END
   END n_88555

   PIN n_88572
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.098 59.997 74.126 60.16 ;
      END
   END n_88572

   PIN n_88589
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.914 59.997 92.942 60.16 ;
      END
   END n_88589

   PIN n_88594
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.938 59.997 77.966 60.16 ;
      END
   END n_88594

   PIN n_88626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 50.226 106.624 50.254 ;
      END
   END n_88626

   PIN n_88646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 42.098 106.624 42.126 ;
      END
   END n_88646

   PIN n_88652
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.962 59.997 78.99 60.16 ;
      END
   END n_88652

   PIN n_88668
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.778 106.624 49.806 ;
      END
   END n_88668

   PIN n_88683
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.85 59.997 92.878 60.16 ;
      END
   END n_88683

   PIN n_88697
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.778 59.997 81.806 60.16 ;
      END
   END n_88697

   PIN n_88703
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.098 59.997 98.126 60.16 ;
      END
   END n_88703

   PIN n_88704
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.714 59.997 81.742 60.16 ;
      END
   END n_88704

   PIN n_88705
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.33 59.997 89.358 60.16 ;
      END
   END n_88705

   PIN n_88706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.874 59.997 77.902 60.16 ;
      END
   END n_88706

   PIN n_88707
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.266 59.997 89.294 60.16 ;
      END
   END n_88707

   PIN n_88708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.202 59.997 89.23 60.16 ;
      END
   END n_88708

   PIN n_88786
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.514 59.997 86.542 60.16 ;
      END
   END n_88786

   PIN n_88805
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.33 59.997 89.358 60.16 ;
      END
   END n_88805

   PIN n_88833
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.922 106.624 39.95 ;
      END
   END n_88833

   PIN n_88835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.49 59.997 85.518 60.16 ;
      END
   END n_88835

   PIN n_88854
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 40.626 106.624 40.654 ;
      END
   END n_88854

   PIN n_89083
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.426 59.997 85.454 60.16 ;
      END
   END n_89083

   PIN n_89164
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.362 59.997 85.39 60.16 ;
      END
   END n_89164

   PIN n_89232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.954 59.997 99.982 60.16 ;
      END
   END n_89232

   PIN n_89272
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.402 59.997 100.43 60.16 ;
      END
   END n_89272

   PIN n_89334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.298 59.997 101.326 60.16 ;
      END
   END n_89334

   PIN n_89338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.018 59.997 100.046 60.16 ;
      END
   END n_89338

   PIN n_89339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.49 59.997 101.518 60.16 ;
      END
   END n_89339

   PIN n_89351
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.186 59.997 99.214 60.16 ;
      END
   END n_89351

   PIN n_89410
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.738 60.078 98.766 60.16 ;
      END
   END n_89410

   PIN n_89426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.634 59.997 99.662 60.16 ;
      END
   END n_89426

   PIN n_89435
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.314 59.997 99.342 60.16 ;
      END
   END n_89435

   PIN n_89436
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.13 59.997 94.158 60.16 ;
      END
   END n_89436

   PIN n_89496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.082 59.997 100.11 60.16 ;
      END
   END n_89496

   PIN n_89517
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.698 59.997 99.726 60.16 ;
      END
   END n_89517

   PIN n_89518
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.058 59.997 99.086 60.16 ;
      END
   END n_89518

   PIN n_89528
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.874 59.997 101.902 60.16 ;
      END
   END n_89528

   PIN n_89581
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.25 59.997 99.278 60.16 ;
      END
   END n_89581

   PIN n_89657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.058 59.997 99.086 60.16 ;
      END
   END n_89657

   PIN n_89673
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.658 59.997 100.686 60.16 ;
      END
   END n_89673

   PIN n_89840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.226 59.997 98.254 60.16 ;
      END
   END n_89840

   PIN n_89892
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.858 106.624 47.886 ;
      END
   END n_89892

   PIN n_89963
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.634 59.997 99.662 60.16 ;
      END
   END n_89963

   PIN n_90020
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 44.85 106.624 44.878 ;
      END
   END n_90020

   PIN n_90052
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.57 59.997 99.598 60.16 ;
      END
   END n_90052

   PIN n_90172
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.682 59.997 93.71 60.16 ;
      END
   END n_90172

   PIN n_90334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.034 59.997 74.062 60.16 ;
      END
   END n_90334

   PIN n_90504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.29 59.997 98.318 60.16 ;
      END
   END n_90504

   PIN n_90645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.082 59.997 100.11 60.16 ;
      END
   END n_90645

   PIN n_90656
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.738 59.997 66.766 60.16 ;
      END
   END n_90656

   PIN n_90669
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.346 106.624 47.374 ;
      END
   END n_90669

   PIN n_90684
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.282 106.624 47.31 ;
      END
   END n_90684

   PIN n_90710
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.45 59.997 86.478 60.16 ;
      END
   END n_90710

   PIN n_90712
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 46.706 106.624 46.734 ;
      END
   END n_90712

   PIN u2_L2_reg_17__Q
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.394 106.624 41.422 ;
      END
   END u2_L2_reg_17__Q

   PIN u2_L2_reg_9__Q
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 40.69 106.624 40.718 ;
      END
   END u2_L2_reg_9__Q

   PIN u2_L3_reg_17__Q
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 45.042 106.624 45.07 ;
      END
   END u2_L3_reg_17__Q

   PIN u2_L3_reg_9__Q
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.93 59.997 98.958 60.16 ;
      END
   END u2_L3_reg_9__Q

   PIN u2_L4_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 35.442 106.624 35.47 ;
      END
   END u2_L4_12_

   PIN u2_L4_19_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.97 59.997 73.998 60.16 ;
      END
   END u2_L4_19_

   PIN u2_L4_22_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.938 59.997 101.966 60.16 ;
      END
   END u2_L4_22_

   PIN u2_L4_29_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 34.162 106.624 34.19 ;
      END
   END u2_L4_29_

   PIN u2_L4_reg_7__Q
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 32.946 106.624 32.974 ;
      END
   END u2_L4_reg_7__Q

   PIN u2_R2_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 39.538 106.624 39.566 ;
      END
   END u2_R2_13_

   PIN u2_R2_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 43.762 106.624 43.79 ;
      END
   END u2_R2_14_

   PIN u2_R2_28_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 37.362 106.624 37.39 ;
      END
   END u2_R2_28_

   PIN u2_R2_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.682 106.624 45.71 ;
      END
   END u2_R2_2_

   PIN u2_R3_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 42.93 106.624 42.958 ;
      END
   END u2_R3_11_

   PIN u2_R3_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.33 106.624 41.358 ;
      END
   END u2_R3_12_

   PIN u2_R3_17_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.266 106.624 41.294 ;
      END
   END u2_R3_17_

   PIN u2_R3_18_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 43.314 106.624 43.342 ;
      END
   END u2_R3_18_

   PIN u2_R3_22_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 49.714 106.624 49.742 ;
      END
   END u2_R3_22_

   PIN u2_R3_23_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 41.97 106.624 41.998 ;
      END
   END u2_R3_23_

   PIN u2_R3_26_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.586 0.0 97.614 0.163 ;
      END
   END u2_R3_26_

   PIN u2_R3_28_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 43.378 106.624 43.406 ;
      END
   END u2_R3_28_

   PIN u2_R3_31_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 45.042 106.624 45.07 ;
      END
   END u2_R3_31_

   PIN u2_R3_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.418 59.997 98.446 60.16 ;
      END
   END u2_R3_3_

   PIN u2_R3_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.906 106.624 41.934 ;
      END
   END u2_R3_4_

   PIN u2_R3_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.09 59.997 103.118 60.16 ;
      END
   END u2_R3_5_

   PIN u2_R3_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 41.65 106.624 41.678 ;
      END
   END u2_R3_8_

   PIN u2_R4_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 106.461 47.794 106.624 47.822 ;
      END
   END u2_R4_10_

   PIN u2_R4_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 44.786 106.624 44.814 ;
      END
   END u2_R4_12_

   PIN u2_R4_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.386 59.997 102.414 60.16 ;
      END
   END u2_R4_14_

   PIN u2_R4_24_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.642 59.997 78.67 60.16 ;
      END
   END u2_R4_24_

   PIN u2_R4_26_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.514 59.997 102.542 60.16 ;
      END
   END u2_R4_26_

   PIN u2_R4_30_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.49 59.997 101.518 60.16 ;
      END
   END u2_R4_30_

   PIN u2_R4_31_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 106.461 41.906 106.624 41.934 ;
      END
   END u2_R4_31_

   PIN u2_uk_K_r_420
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.13 59.997 102.158 60.16 ;
      END
   END u2_uk_K_r_420

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 106.624 60.16 ;
      LAYER V1 ;
         RECT 0.0 0.0 106.624 60.16 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 106.624 60.16 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 106.624 60.16 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 106.624 60.16 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 106.624 60.16 ;
      LAYER M1 ;
         RECT 0.0 0.0 106.624 60.16 ;
   END
END h1_mgc_des_perf_a

MACRO h0_mgc_des_perf_a
   CLASS BLOCK ;
   FOREIGN h0 ;
   ORIGIN 0 0 ;
   SIZE 89.6 BY 94.979 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN2124_n_92148
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 43.25 89.6 43.278 ;
      END
   END FE_OFN2124_n_92148

   PIN FE_OFN2215_n_2854
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.322 0.0 38.35 0.163 ;
      END
   END FE_OFN2215_n_2854

   PIN g202734_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 47.346 89.6 47.374 ;
      END
   END g202734_p

   PIN g289278_p2
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.362 0.0 29.39 0.163 ;
      END
   END g289278_p2

   PIN g289637_p1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.306 0.0 48.334 0.163 ;
      END
   END g289637_p1

   PIN g291339_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.226 0.0 42.254 0.163 ;
      END
   END g291339_p

   PIN g301491_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.658 0.163 12.686 ;
      END
   END g301491_p

   PIN g302166_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.706 0.163 22.734 ;
      END
   END g302166_p

   PIN key_c_r_26__2568
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.89 0.0 27.918 0.163 ;
      END
   END key_c_r_26__2568

   PIN n_10300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.978 0.0 37.006 0.163 ;
      END
   END n_10300

   PIN n_10543
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.21 0.0 44.238 0.163 ;
      END
   END n_10543

   PIN n_10664
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.106 0.0 45.134 0.163 ;
      END
   END n_10664

   PIN n_11092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.722 0.0 44.75 0.163 ;
      END
   END n_11092

   PIN n_11160
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.298 0.0 37.326 0.163 ;
      END
   END n_11160

   PIN n_11190
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.522 0.0 41.55 0.163 ;
      END
   END n_11190

   PIN n_11283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.042 0.0 37.07 0.163 ;
      END
   END n_11283

   PIN n_116769
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.858 0.0 63.886 0.163 ;
      END
   END n_116769

   PIN n_116784
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.45 0.0 6.478 0.163 ;
      END
   END n_116784

   PIN n_117640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.362 0.0 45.39 0.163 ;
      END
   END n_117640

   PIN n_117987
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.362 0.0 61.39 0.163 ;
      END
   END n_117987

   PIN n_1204
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.818 0.0 64.846 0.163 ;
      END
   END n_1204

   PIN n_1209
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.026 0.163 55.054 ;
      END
   END n_1209

   PIN n_12805
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 0.0 25.614 0.163 ;
      END
   END n_12805

   PIN n_12937
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.706 0.0 30.734 0.163 ;
      END
   END n_12937

   PIN n_12977
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.522 0.0 25.55 0.163 ;
      END
   END n_12977

   PIN n_1417
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.762 0.0 59.79 0.163 ;
      END
   END n_1417

   PIN n_14736
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.306 0.0 72.334 0.163 ;
      END
   END n_14736

   PIN n_1579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.842 0.0 65.87 0.163 ;
      END
   END n_1579

   PIN n_17638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.074 0.0 73.102 0.163 ;
      END
   END n_17638

   PIN n_18022
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.026 0.0 87.054 0.163 ;
      END
   END n_18022

   PIN n_18160
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.914 89.6 4.942 ;
      END
   END n_18160

   PIN n_2208
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.01 0.163 9.038 ;
      END
   END n_2208

   PIN n_2598
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.626 0.163 16.654 ;
      END
   END n_2598

   PIN n_3390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.626 0.163 16.654 ;
      END
   END n_3390

   PIN n_3453
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.722 0.163 12.75 ;
      END
   END n_3453

   PIN n_3518
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.426 0.0 29.454 0.163 ;
      END
   END n_3518

   PIN n_3653
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.85 0.163 12.878 ;
      END
   END n_3653

   PIN n_3919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.482 0.163 26.51 ;
      END
   END n_3919

   PIN n_4023
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.682 0.0 21.71 0.163 ;
      END
   END n_4023

   PIN n_4025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.402 0.163 20.43 ;
      END
   END n_4025

   PIN n_4166
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.746 0.0 21.774 0.163 ;
      END
   END n_4166

   PIN n_4717
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.466 0.163 20.494 ;
      END
   END n_4717

   PIN n_4718
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.818 0.163 16.846 ;
      END
   END n_4718

   PIN n_4927
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.69 0.163 16.718 ;
      END
   END n_4927

   PIN n_5717
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.826 0.163 35.854 ;
      END
   END n_5717

   PIN n_66187
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 20.466 89.6 20.494 ;
      END
   END n_66187

   PIN n_66261
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 20.53 89.6 20.558 ;
      END
   END n_66261

   PIN n_7078
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.57 0.0 75.598 0.163 ;
      END
   END n_7078

   PIN n_7087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 46.002 0.0 46.03 0.163 ;
      END
   END n_7087

   PIN n_7431
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.634 0.0 67.662 0.163 ;
      END
   END n_7431

   PIN n_7877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.802 0.0 50.83 0.163 ;
      END
   END n_7877

   PIN n_8063
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.978 0.0 45.006 0.163 ;
      END
   END n_8063

   PIN n_8726
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 49.97 0.0 49.998 0.163 ;
      END
   END n_8726

   PIN n_8829
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.418 0.0 50.446 0.163 ;
      END
   END n_8829

   PIN n_91001
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 39.602 89.6 39.63 ;
      END
   END n_91001

   PIN n_9103
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.522 0.0 49.55 0.163 ;
      END
   END n_9103

   PIN n_91121
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 28.082 89.6 28.11 ;
      END
   END n_91121

   PIN n_91266
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 8.946 89.6 8.974 ;
      END
   END n_91266

   PIN n_91489
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 9.138 89.6 9.166 ;
      END
   END n_91489

   PIN n_91525
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 32.05 89.6 32.078 ;
      END
   END n_91525

   PIN n_91573
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.978 89.6 5.006 ;
      END
   END n_91573

   PIN n_91692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 31.858 89.6 31.886 ;
      END
   END n_91692

   PIN n_91814
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 32.114 89.6 32.142 ;
      END
   END n_91814

   PIN n_91815
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.338 89.6 4.366 ;
      END
   END n_91815

   PIN n_91824
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 39.73 89.6 39.758 ;
      END
   END n_91824

   PIN n_91825
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 43.442 89.6 43.47 ;
      END
   END n_91825

   PIN n_91826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 31.922 89.6 31.95 ;
      END
   END n_91826

   PIN n_91828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 35.826 89.6 35.854 ;
      END
   END n_91828

   PIN n_91839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 35.89 89.6 35.918 ;
      END
   END n_91839

   PIN n_91845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 9.01 89.6 9.038 ;
      END
   END n_91845

   PIN n_92019
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 8.882 89.6 8.91 ;
      END
   END n_92019

   PIN n_92117
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 35.954 89.6 35.982 ;
      END
   END n_92117

   PIN n_92305
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 5.042 89.6 5.07 ;
      END
   END n_92305

   PIN n_92419
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 36.018 89.6 36.046 ;
      END
   END n_92419

   PIN n_92502
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 89.437 3.698 89.6 3.726 ;
      END
   END n_92502

   PIN n_92510
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 9.074 89.6 9.102 ;
      END
   END n_92510

   PIN n_92511
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 43.506 89.6 43.534 ;
      END
   END n_92511

   PIN n_9282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.058 0.0 51.086 0.163 ;
      END
   END n_9282

   PIN n_95488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 47.41 89.6 47.438 ;
      END
   END n_95488

   PIN n_95562
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 5.106 89.6 5.134 ;
      END
   END n_95562

   PIN n_95579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 3.826 89.6 3.854 ;
      END
   END n_95579

   PIN n_95580
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 47.474 89.6 47.502 ;
      END
   END n_95580

   PIN n_95719
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 51.186 89.6 51.214 ;
      END
   END n_95719

   PIN n_95756
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 9.202 89.6 9.23 ;
      END
   END n_95756

   PIN n_95826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.518 3.506 89.6 3.534 ;
      END
   END n_95826

   PIN n_95913
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 55.026 89.6 55.054 ;
      END
   END n_95913

   PIN n_95976
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 9.266 89.6 9.294 ;
      END
   END n_95976

   PIN n_96109
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 47.538 89.6 47.566 ;
      END
   END n_96109

   PIN n_96227
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 51.25 89.6 51.278 ;
      END
   END n_96227

   PIN n_96448
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 9.33 89.6 9.358 ;
      END
   END n_96448

   PIN n_96488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 12.786 89.6 12.814 ;
      END
   END n_96488

   PIN n_9734
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.098 0.0 50.126 0.163 ;
      END
   END n_9734

   PIN u0_L0_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.674 0.0 2.702 0.163 ;
      END
   END u0_L0_10_

   PIN u0_L0_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.65 0.0 25.678 0.163 ;
      END
   END u0_L0_4_

   PIN u0_L0_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.786 0.0 44.814 0.163 ;
      END
   END u0_L0_6_

   PIN u0_L1_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.394 0.0 73.422 0.163 ;
      END
   END u0_L1_10_

   PIN u0_L1_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.242 0.0 56.27 0.163 ;
      END
   END u0_L1_1_

   PIN u0_R0_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.866 0.0 34.894 0.163 ;
      END
   END u0_R0_23_

   PIN u0_R0_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.058 0.0 59.086 0.163 ;
      END
   END u0_R0_28_

   PIN u1_key_r_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 42.61 89.6 42.638 ;
      END
   END u1_key_r_28_

   PIN FE_OFN1268_n_3950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.402 0.163 28.43 ;
      END
   END FE_OFN1268_n_3950

   PIN FE_OFN1270_n_6370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.986 0.163 32.014 ;
      END
   END FE_OFN1270_n_6370

   PIN FE_OFN1342_n_5733
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.506 0.0 35.534 0.163 ;
      END
   END FE_OFN1342_n_5733

   PIN FE_OFN1346_n_1012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.146 0.0 60.174 0.163 ;
      END
   END FE_OFN1346_n_1012

   PIN FE_OFN1882_n_1371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.802 0.163 26.83 ;
      END
   END FE_OFN1882_n_1371

   PIN FE_OFN2123_n_92148
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 28.21 89.6 28.238 ;
      END
   END FE_OFN2123_n_92148

   PIN FE_OFN2356_n_1288
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.514 0.0 46.542 0.163 ;
      END
   END FE_OFN2356_n_1288

   PIN FE_OFN749_n_15670
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.922 0.0 63.95 0.163 ;
      END
   END FE_OFN749_n_15670

   PIN desIn_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.106 0.163 5.134 ;
      END
   END desIn_13_

   PIN desIn_31_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.042 0.163 5.07 ;
      END
   END desIn_31_

   PIN desIn_38_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.026 94.815 87.054 94.978 ;
      END
   END desIn_38_

   PIN desIn_50_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.786 0.163 12.814 ;
      END
   END desIn_50_

   PIN g303844_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.346 0.0 79.374 0.163 ;
      END
   END g303844_db

   PIN g303844_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.186 0.0 83.214 0.163 ;
      END
   END g303844_sb

   PIN g321474_db
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.61 0.0 2.638 0.163 ;
      END
   END g321474_db

   PIN g321474_sb
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.642 0.0 22.67 0.163 ;
      END
   END g321474_sb

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.518 42.482 89.6 42.51 ;
      END
   END ispd_clk

   PIN key_b_r_16__28_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 94.815 25.614 94.978 ;
      END
   END key_b_r_16__28_

   PIN key_c_r_25__2513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.21 94.815 28.238 94.978 ;
      END
   END key_c_r_25__2513

   PIN n_10016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.202 0.0 33.23 0.163 ;
      END
   END n_10016

   PIN n_10047
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.234 0.0 37.262 0.163 ;
      END
   END n_10047

   PIN n_10087
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.33 0.0 41.358 0.163 ;
      END
   END n_10087

   PIN n_10299
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.338 0.0 44.366 0.163 ;
      END
   END n_10299

   PIN n_10307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.266 0.0 33.294 0.163 ;
      END
   END n_10307

   PIN n_10322
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.946 0.0 40.974 0.163 ;
      END
   END n_10322

   PIN n_10332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.17 0.0 37.198 0.082 ;
      END
   END n_10332

   PIN n_10534
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.546 0.0 42.574 0.163 ;
      END
   END n_10534

   PIN n_10560
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.138 0.0 33.166 0.163 ;
      END
   END n_10560

   PIN n_10579
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.434 0.0 48.462 0.163 ;
      END
   END n_10579

   PIN n_10628
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.394 0.0 41.422 0.082 ;
      END
   END n_10628

   PIN n_10707
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.034 0.0 50.062 0.163 ;
      END
   END n_10707

   PIN n_10905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.314 0.0 43.342 0.163 ;
      END
   END n_10905

   PIN n_116767
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.81 0.0 69.838 0.163 ;
      END
   END n_116767

   PIN n_116774
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.138 0.0 73.166 0.163 ;
      END
   END n_116774

   PIN n_117986
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.514 0.0 62.542 0.163 ;
      END
   END n_117986

   PIN n_11904
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.098 0.0 42.126 0.163 ;
      END
   END n_11904

   PIN n_11922
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.298 0.0 45.326 0.163 ;
      END
   END n_11922

   PIN n_12137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.914 0.0 36.942 0.163 ;
      END
   END n_12137

   PIN n_1241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.49 0.0 29.518 0.163 ;
      END
   END n_1241

   PIN n_12565
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.298 0.0 29.326 0.163 ;
      END
   END n_12565

   PIN n_1323
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.61 0.0 74.638 0.163 ;
      END
   END n_1323

   PIN n_14285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.37 0.0 72.398 0.163 ;
      END
   END n_14285

   PIN n_15830
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.306 0.0 56.334 0.163 ;
      END
   END n_15830

   PIN n_15918
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.306 0.0 56.334 0.163 ;
      END
   END n_15918

   PIN n_16285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.658 0.0 68.686 0.163 ;
      END
   END n_16285

   PIN n_16293
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.082 0.0 60.11 0.082 ;
      END
   END n_16293

   PIN n_16596
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.514 0.0 70.542 0.163 ;
      END
   END n_16596

   PIN n_16597
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.09 0.0 71.118 0.163 ;
      END
   END n_16597

   PIN n_16611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.922 0.0 63.95 0.163 ;
      END
   END n_16611

   PIN n_1662
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.626 0.163 24.654 ;
      END
   END n_1662

   PIN n_16731
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.018 0.0 60.046 0.163 ;
      END
   END n_16731

   PIN n_16854
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.938 0.0 69.966 0.163 ;
      END
   END n_16854

   PIN n_1686
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.562 0.163 24.59 ;
      END
   END n_1686

   PIN n_16882
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.018 0.0 60.046 0.163 ;
      END
   END n_16882

   PIN n_17069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.962 0.0 70.99 0.163 ;
      END
   END n_17069

   PIN n_17155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.106 0.0 69.134 0.163 ;
      END
   END n_17155

   PIN n_1844
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.922 0.163 23.95 ;
      END
   END n_1844

   PIN n_1916
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.546 0.0 2.574 0.163 ;
      END
   END n_1916

   PIN n_2108
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.642 0.163 22.67 ;
      END
   END n_2108

   PIN n_2210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.514 0.0 6.542 0.163 ;
      END
   END n_2210

   PIN n_2597
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.906 0.0 17.934 0.163 ;
      END
   END n_2597

   PIN n_2610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.546 0.0 2.574 0.163 ;
      END
   END n_2610

   PIN n_2611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.25 0.0 83.278 0.163 ;
      END
   END n_2611

   PIN n_2721
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.946 0.163 8.974 ;
      END
   END n_2721

   PIN n_2854
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.226 0.0 10.254 0.163 ;
      END
   END n_2854

   PIN n_2883
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.562 0.163 16.59 ;
      END
   END n_2883

   PIN n_2885
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.73 0.082 23.758 ;
      END
   END n_2885

   PIN n_3058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.386 0.0 6.414 0.163 ;
      END
   END n_3058

   PIN n_3098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.498 0.163 16.526 ;
      END
   END n_3098

   PIN n_3175
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.53 0.163 20.558 ;
      END
   END n_3175

   PIN n_3238
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.754 0.163 16.782 ;
      END
   END n_3238

   PIN n_3397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.69 0.163 24.718 ;
      END
   END n_3397

   PIN n_3431
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.466 0.163 20.494 ;
      END
   END n_3431

   PIN n_3517
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.786 0.163 12.814 ;
      END
   END n_3517

   PIN n_3652
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.434 0.163 16.462 ;
      END
   END n_3652

   PIN n_3798
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.466 0.163 28.494 ;
      END
   END n_3798

   PIN n_3856
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.882 0.163 8.91 ;
      END
   END n_3856

   PIN n_3942
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.842 0.163 25.87 ;
      END
   END n_3942

   PIN n_3949
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.922 0.163 31.95 ;
      END
   END n_3949

   PIN n_4410
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.37 0.163 16.398 ;
      END
   END n_4410

   PIN n_4867
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.05 0.163 32.078 ;
      END
   END n_4867

   PIN n_4868
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.386 0.0 6.414 0.163 ;
      END
   END n_4868

   PIN n_4933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.618 0.0 21.646 0.163 ;
      END
   END n_4933

   PIN n_5261
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.762 0.163 27.79 ;
      END
   END n_5261

   PIN n_5296
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.402 0.163 20.43 ;
      END
   END n_5296

   PIN n_65597
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.85 89.6 4.878 ;
      END
   END n_65597

   PIN n_65740
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 16.626 89.6 16.654 ;
      END
   END n_65740

   PIN n_65860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 20.402 89.6 20.43 ;
      END
   END n_65860

   PIN n_6598
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.026 0.0 63.054 0.163 ;
      END
   END n_6598

   PIN n_66080
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.518 4.21 89.6 4.238 ;
      END
   END n_66080

   PIN n_66260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 24.242 89.6 24.27 ;
      END
   END n_66260

   PIN n_6675
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.466 0.0 52.494 0.163 ;
      END
   END n_6675

   PIN n_7855
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.402 0.0 52.43 0.163 ;
      END
   END n_7855

   PIN n_8357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.122 0.0 51.15 0.163 ;
      END
   END n_8357

   PIN n_8586
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.738 0.0 50.766 0.163 ;
      END
   END n_8586

   PIN n_8587
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.034 0.0 50.062 0.163 ;
      END
   END n_8587

   PIN n_8743
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.85 0.0 36.878 0.163 ;
      END
   END n_8743

   PIN n_8902
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.906 0.0 41.934 0.163 ;
      END
   END n_8902

   PIN n_91003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 35.57 89.6 35.598 ;
      END
   END n_91003

   PIN n_91051
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 89.518 3.506 89.6 3.534 ;
      END
   END n_91051

   PIN n_91073
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.578 0.0 86.606 0.163 ;
      END
   END n_91073

   PIN n_91091
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 31.986 89.6 32.014 ;
      END
   END n_91091

   PIN n_91165
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.082 89.6 4.11 ;
      END
   END n_91165

   PIN n_91268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.09 0.0 87.118 0.163 ;
      END
   END n_91268

   PIN n_91345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.786 89.6 4.814 ;
      END
   END n_91345

   PIN n_91373
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.858 0.0 87.886 0.163 ;
      END
   END n_91373

   PIN n_91534
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 28.018 89.6 28.046 ;
      END
   END n_91534

   PIN n_91579
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.018 89.6 4.046 ;
      END
   END n_91579

   PIN n_92127
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 35.762 89.6 35.79 ;
      END
   END n_92127

   PIN n_92142
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 35.698 89.6 35.726 ;
      END
   END n_92142

   PIN n_92144
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 39.666 89.6 39.694 ;
      END
   END n_92144

   PIN n_92271
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 28.146 89.6 28.174 ;
      END
   END n_92271

   PIN n_92319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.722 89.6 4.75 ;
      END
   END n_92319

   PIN n_92482
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 35.634 89.6 35.662 ;
      END
   END n_92482

   PIN n_934
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.074 0.0 65.102 0.163 ;
      END
   END n_934

   PIN n_935
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.098 0.0 34.126 0.163 ;
      END
   END n_935

   PIN n_9426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.786 0.0 36.814 0.163 ;
      END
   END n_9426

   PIN n_9428
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.714 0.0 49.742 0.163 ;
      END
   END n_9428

   PIN n_9499
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.17 0.0 37.198 0.163 ;
      END
   END n_9499

   PIN n_95152
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 47.154 89.6 47.182 ;
      END
   END n_95152

   PIN n_95239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 43.378 89.6 43.406 ;
      END
   END n_95239

   PIN n_95318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 43.314 89.6 43.342 ;
      END
   END n_95318

   PIN n_95323
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.658 89.6 4.686 ;
      END
   END n_95323

   PIN n_95363
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 3.762 89.6 3.79 ;
      END
   END n_95363

   PIN n_95397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.594 89.6 4.622 ;
      END
   END n_95397

   PIN n_95412
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.53 89.6 4.558 ;
      END
   END n_95412

   PIN n_95416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.466 89.6 4.494 ;
      END
   END n_95416

   PIN n_95587
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 4.402 89.6 4.43 ;
      END
   END n_95587

   PIN n_95604
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.518 3.634 89.6 3.662 ;
      END
   END n_95604

   PIN n_95698
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 47.218 89.6 47.246 ;
      END
   END n_95698

   PIN n_95810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 47.282 89.6 47.31 ;
      END
   END n_95810

   PIN n_96003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 51.122 89.6 51.15 ;
      END
   END n_96003

   PIN n_96004
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 3.954 89.6 3.982 ;
      END
   END n_96004

   PIN n_96232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 89.437 3.89 89.6 3.918 ;
      END
   END n_96232

   PIN n_96447
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 89.437 3.634 89.6 3.662 ;
      END
   END n_96447

   PIN n_9741
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.106 0.0 37.134 0.163 ;
      END
   END n_9741

   PIN n_9764
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.786 0.0 44.814 0.163 ;
      END
   END n_9764

   PIN u0_IP_64__1294
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.018 0.0 68.046 0.163 ;
      END
   END u0_IP_64__1294

   PIN u0_R0_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.162 0.0 74.19 0.163 ;
      END
   END u0_R0_10_

   PIN u0_R0_20_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.162 0.0 66.19 0.163 ;
      END
   END u0_R0_20_

   PIN u0_R0_24_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.194 0.0 46.222 0.163 ;
      END
   END u0_R0_24_

   PIN u0_R0_26_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.81 0.0 61.838 0.163 ;
      END
   END u0_R0_26_

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 89.6 94.979 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 89.6 94.979 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 89.6 94.979 ;
      LAYER V1 ;
         RECT 0.0 0.0 89.6 94.979 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 89.6 94.979 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 89.6 94.979 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 89.6 94.979 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 89.6 94.979 ;
      LAYER M1 ;
         RECT 0.0 0.0 89.6 94.979 ;
   END
END h0_mgc_des_perf_a

MACRO h4_mgc_edit_dist_a
   CLASS BLOCK ;
   FOREIGN h4 ;
   ORIGIN 0 0 ;
   SIZE 53.376 BY 76.8 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN57649_FE_OFN47241_n_6273_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.482 0.163 42.51 ;
      END
   END FE_OCPN57649_FE_OFN47241_n_6273_bar

   PIN FE_OCPN61274_n_33700_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 5.426 53.376 5.454 ;
      END
   END FE_OCPN61274_n_33700_bar

   PIN FE_OCPN61430_n_31308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.57 0.163 75.598 ;
      END
   END FE_OCPN61430_n_31308

   PIN FE_OCPN61542_FE_OFN47238_mux_k_ln251_z_5__4323813_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.322 0.163 46.35 ;
      END
   END FE_OCPN61542_FE_OFN47238_mux_k_ln251_z_5__4323813_bar

   PIN FE_OCPN61544_n_35219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.514 0.163 38.542 ;
      END
   END FE_OCPN61544_n_35219

   PIN FE_OCPN61546_n_35219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 23.154 0.082 23.182 ;
      END
   END FE_OCPN61546_n_35219

   PIN FE_OCPN62339_n_65283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.762 0.163 51.79 ;
      END
   END FE_OCPN62339_n_65283

   PIN FE_OCPN63165_n_34645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.242 0.163 24.27 ;
      END
   END FE_OCPN63165_n_34645

   PIN FE_OCPN63166_n_34645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 21.106 0.163 21.134 ;
      END
   END FE_OCPN63166_n_34645

   PIN FE_OCPN63167_n_34645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.026 0.163 31.054 ;
      END
   END FE_OCPN63167_n_34645

   PIN FE_OCPN63170_n_34645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.922 0.163 23.95 ;
      END
   END FE_OCPN63170_n_34645

   PIN FE_OCPN63172_n_34609
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.666 0.163 15.694 ;
      END
   END FE_OCPN63172_n_34609

   PIN FE_OCPN63184_n_34610
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.994 0.163 35.022 ;
      END
   END FE_OCPN63184_n_34610

   PIN FE_OCPN63185_n_34610
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.002 0.163 22.03 ;
      END
   END FE_OCPN63185_n_34610

   PIN FE_OCPN63189_FE_OFN47238_mux_k_ln251_z_5__4323813_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.778 0.163 25.806 ;
      END
   END FE_OCPN63189_FE_OFN47238_mux_k_ln251_z_5__4323813_bar

   PIN FE_OCPN63285_n_35466
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.61 0.163 34.638 ;
      END
   END FE_OCPN63285_n_35466

   PIN FE_OCPN63376_FE_OFN38554_n_42605
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.274 0.163 60.302 ;
      END
   END FE_OCPN63376_FE_OFN38554_n_42605

   PIN FE_OCPN63733_n_34650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 22.002 0.163 22.03 ;
      END
   END FE_OCPN63733_n_34650

   PIN FE_OCPN63744_n_34677
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.882 0.163 32.91 ;
      END
   END FE_OCPN63744_n_34677

   PIN FE_OFN27591_n_36720
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 66.354 0.163 66.382 ;
      END
   END FE_OFN27591_n_36720

   PIN FE_OFN27671_n_36750
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 71.282 0.163 71.31 ;
      END
   END FE_OFN27671_n_36750

   PIN FE_OFN27677_n_36830
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.114 0.163 72.142 ;
      END
   END FE_OFN27677_n_36830

   PIN FE_OFN27695_n_36869
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 43.954 53.376 43.982 ;
      END
   END FE_OFN27695_n_36869

   PIN FE_OFN27737_n_36719
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.722 0.163 68.75 ;
      END
   END FE_OFN27737_n_36719

   PIN FE_OFN27793_n_36739
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.306 0.163 72.334 ;
      END
   END FE_OFN27793_n_36739

   PIN FE_OFN27858_n_36176
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.634 0.163 75.662 ;
      END
   END FE_OFN27858_n_36176

   PIN FE_OFN27943_n_36631
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.826 0.0 35.854 0.163 ;
      END
   END FE_OFN27943_n_36631

   PIN FE_OFN27945_n_36632
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.378 0.0 35.406 0.163 ;
      END
   END FE_OFN27945_n_36632

   PIN FE_OFN28066_n_36155
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.866 0.0 34.894 0.163 ;
      END
   END FE_OFN28066_n_36155

   PIN FE_OFN28109_n_36231
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.73 53.376 31.758 ;
      END
   END FE_OFN28109_n_36231

   PIN FE_OFN28150_n_36991
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 54.642 53.376 54.67 ;
      END
   END FE_OFN28150_n_36991

   PIN FE_OFN28264_n_36480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 48.882 53.376 48.91 ;
      END
   END FE_OFN28264_n_36480

   PIN FE_OFN30064_n_39931
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 28.914 53.376 28.942 ;
      END
   END FE_OFN30064_n_39931

   PIN FE_OFN32324_g2_n_3744391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 48.498 53.376 48.526 ;
      END
   END FE_OFN32324_g2_n_3744391

   PIN FE_OFN32385_n_21110
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 43.186 53.376 43.214 ;
      END
   END FE_OFN32385_n_21110

   PIN FE_OFN32386_n_21110
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 52.466 0.163 52.494 ;
      END
   END FE_OFN32386_n_21110

   PIN FE_OFN32390_n_59356
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.442 0.082 51.47 ;
      END
   END FE_OFN32390_n_59356

   PIN FE_OFN34192_n_82
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 44.402 53.376 44.43 ;
      END
   END FE_OFN34192_n_82

   PIN FE_OFN34385_n_7916
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.914 0.163 68.942 ;
      END
   END FE_OFN34385_n_7916

   PIN FE_OFN35296_n_5226969_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 30.45 53.376 30.478 ;
      END
   END FE_OFN35296_n_5226969_bar

   PIN FE_OFN35387_eq_15876_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 39.282 0.163 39.31 ;
      END
   END FE_OFN35387_eq_15876_46_n_18

   PIN FE_OFN35405_eq_15784_44_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.778 76.637 17.806 76.8 ;
      END
   END FE_OFN35405_eq_15784_44_n_18

   PIN FE_OFN35416_eq_15782_44_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.386 76.637 6.414 76.8 ;
      END
   END FE_OFN35416_eq_15782_44_n_18

   PIN FE_OFN35557_n_48868
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.346 0.163 55.374 ;
      END
   END FE_OFN35557_n_48868

   PIN FE_OFN35566_n_48307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.938 0.163 45.966 ;
      END
   END FE_OFN35566_n_48307

   PIN FE_OFN35724_n_49478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.13 76.637 6.158 76.8 ;
      END
   END FE_OFN35724_n_49478

   PIN FE_OFN35827_n_43179
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.402 0.163 12.43 ;
      END
   END FE_OFN35827_n_43179

   PIN FE_OFN35833_n_41388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.682 0.163 5.71 ;
      END
   END FE_OFN35833_n_41388

   PIN FE_OFN35980_n_51064
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.546 0.163 58.574 ;
      END
   END FE_OFN35980_n_51064

   PIN FE_OFN35982_n_51575
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.842 0.163 57.87 ;
      END
   END FE_OFN35982_n_51575

   PIN FE_OFN36039_n_49324
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.562 0.163 56.59 ;
      END
   END FE_OFN36039_n_49324

   PIN FE_OFN36056_n_43053
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.266 0.0 9.294 0.163 ;
      END
   END FE_OFN36056_n_43053

   PIN FE_OFN36062_n_40128
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.314 0.163 11.342 ;
      END
   END FE_OFN36062_n_40128

   PIN FE_OFN36065_n_48779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.074 0.163 49.102 ;
      END
   END FE_OFN36065_n_48779

   PIN FE_OFN36096_n_48764
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.698 0.0 43.726 0.163 ;
      END
   END FE_OFN36096_n_48764

   PIN FE_OFN36240_n_48902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.37 0.163 48.398 ;
      END
   END FE_OFN36240_n_48902

   PIN FE_OFN36242_n_49413
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.81 0.163 45.838 ;
      END
   END FE_OFN36242_n_49413

   PIN FE_OFN36289_n_35472
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.122 0.163 19.15 ;
      END
   END FE_OFN36289_n_35472

   PIN FE_OFN36290_n_35472
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.138 0.163 17.166 ;
      END
   END FE_OFN36290_n_35472

   PIN FE_OFN36305_sub_ln263_unr88_z_4__4328191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.786 0.163 28.814 ;
      END
   END FE_OFN36305_sub_ln263_unr88_z_4__4328191

   PIN FE_OFN36306_sub_ln263_unr88_z_4__4328191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.85 0.163 28.878 ;
      END
   END FE_OFN36306_sub_ln263_unr88_z_4__4328191

   PIN FE_OFN36312_n_41464
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.858 0.163 31.886 ;
      END
   END FE_OFN36312_n_41464

   PIN FE_OFN36434_n_51052
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.386 76.637 6.414 76.8 ;
      END
   END FE_OFN36434_n_51052

   PIN FE_OFN36478_n_39632
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 46.066 0.163 46.094 ;
      END
   END FE_OFN36478_n_39632

   PIN FE_OFN36488_n_35474
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.226 0.163 18.254 ;
      END
   END FE_OFN36488_n_35474

   PIN FE_OFN36489_n_35474
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.866 0.082 34.894 ;
      END
   END FE_OFN36489_n_35474

   PIN FE_OFN36543_n_49063
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 37.426 0.163 37.454 ;
      END
   END FE_OFN36543_n_49063

   PIN FE_OFN36564_n_48859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.386 0.163 62.414 ;
      END
   END FE_OFN36564_n_48859

   PIN FE_OFN36573_n_48806
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.666 0.0 39.694 0.163 ;
      END
   END FE_OFN36573_n_48806

   PIN FE_OFN36582_n_34613
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.882 0.082 16.91 ;
      END
   END FE_OFN36582_n_34613

   PIN FE_OFN36613_n_49060
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 5.362 0.163 5.39 ;
      END
   END FE_OFN36613_n_49060

   PIN FE_OFN36690_n_34610
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.154 0.163 15.182 ;
      END
   END FE_OFN36690_n_34610

   PIN FE_OFN36698_n_43262
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.21 0.163 20.238 ;
      END
   END FE_OFN36698_n_43262

   PIN FE_OFN36710_n_39974
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.938 0.163 5.966 ;
      END
   END FE_OFN36710_n_39974

   PIN FE_OFN36729_n_35568
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.522 0.163 25.55 ;
      END
   END FE_OFN36729_n_35568

   PIN FE_OFN36733_n_35568
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 21.362 0.163 21.39 ;
      END
   END FE_OFN36733_n_35568

   PIN FE_OFN36770_n_40005
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.49 0.163 5.518 ;
      END
   END FE_OFN36770_n_40005

   PIN FE_OFN36771_n_41490
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.162 0.163 34.19 ;
      END
   END FE_OFN36771_n_41490

   PIN FE_OFN36774_n_39746
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.37 0.163 32.398 ;
      END
   END FE_OFN36774_n_39746

   PIN FE_OFN36787_sub_14956_48_n_104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.01 0.163 9.038 ;
      END
   END FE_OFN36787_sub_14956_48_n_104

   PIN FE_OFN37075_sub_15040_54_n_115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.21 0.163 36.238 ;
      END
   END FE_OFN37075_sub_15040_54_n_115

   PIN FE_OFN37708_n_42708
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 1.906 53.376 1.934 ;
      END
   END FE_OFN37708_n_42708

   PIN FE_OFN38237_sub_15041_54_n_115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.178 0.163 40.206 ;
      END
   END FE_OFN38237_sub_15041_54_n_115

   PIN FE_OFN38498_n_42702
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.002 0.163 46.03 ;
      END
   END FE_OFN38498_n_42702

   PIN FE_OFN38572_n_35480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.002 0.082 14.03 ;
      END
   END FE_OFN38572_n_35480

   PIN FE_OFN41497_sub_15040_54_n_63
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.202 0.163 17.23 ;
      END
   END FE_OFN41497_sub_15040_54_n_63

   PIN FE_OFN41895_n_226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 48.562 53.376 48.59 ;
      END
   END FE_OFN41895_n_226

   PIN FE_OFN41977_n_228
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 47.538 53.376 47.566 ;
      END
   END FE_OFN41977_n_228

   PIN FE_OFN43137_n_35287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.242 0.082 64.27 ;
      END
   END FE_OFN43137_n_35287

   PIN FE_OFN43147_n_35287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 40.818 53.376 40.846 ;
      END
   END FE_OFN43147_n_35287

   PIN FE_OFN44003_n_35331
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 71.282 53.376 71.31 ;
      END
   END FE_OFN44003_n_35331

   PIN FE_OFN46305_n_35331
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 40.69 53.376 40.718 ;
      END
   END FE_OFN46305_n_35331

   PIN FE_OFN46746_n_57645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.474 0.163 63.502 ;
      END
   END FE_OFN46746_n_57645

   PIN FE_OFN46835_n_18055
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 62.962 53.376 62.99 ;
      END
   END FE_OFN46835_n_18055

   PIN FE_OFN46837_n_5223349_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 65.906 53.376 65.934 ;
      END
   END FE_OFN46837_n_5223349_bar

   PIN FE_OFN47466_sub_15040_54_n_63
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.13 0.163 22.158 ;
      END
   END FE_OFN47466_sub_15040_54_n_63

   PIN FE_OFN47467_sub_15040_54_n_63
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.77 0.163 22.798 ;
      END
   END FE_OFN47467_sub_15040_54_n_63

   PIN FE_OFN47469_sub_15027_54_n_55
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.674 0.163 34.702 ;
      END
   END FE_OFN47469_sub_15027_54_n_55

   PIN FE_OFN48512_n_59356
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.026 0.163 23.054 ;
      END
   END FE_OFN48512_n_59356

   PIN FE_OFN49008_n_39642
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.026 0.163 15.054 ;
      END
   END FE_OFN49008_n_39642

   PIN FE_OFN49020_n_42611
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.474 0.163 47.502 ;
      END
   END FE_OFN49020_n_42611

   PIN FE_OFN49964_n_48908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.242 0.163 72.27 ;
      END
   END FE_OFN49964_n_48908

   PIN FE_OFN49999_n_49354
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.41 0.163 55.438 ;
      END
   END FE_OFN49999_n_49354

   PIN FE_OFN50041_n_49465
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.498 0.163 40.526 ;
      END
   END FE_OFN50041_n_49465

   PIN FE_OFN50111_n_49480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 49.074 0.163 49.102 ;
      END
   END FE_OFN50111_n_49480

   PIN FE_OFN50218_n_51418
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.138 0.163 49.166 ;
      END
   END FE_OFN50218_n_51418

   PIN FE_OFN50523_n_57647
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.178 0.163 72.206 ;
      END
   END FE_OFN50523_n_57647

   PIN FE_OFN50623_n_57653
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 47.986 0.163 48.014 ;
      END
   END FE_OFN50623_n_57653

   PIN FE_OFN54179_n_57047
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.426 76.637 29.454 76.8 ;
      END
   END FE_OFN54179_n_57047

   PIN FE_OFN54264_n_57053
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.034 76.637 26.062 76.8 ;
      END
   END FE_OFN54264_n_57053

   PIN FE_OFN70124_n_36963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 75.186 0.163 75.214 ;
      END
   END FE_OFN70124_n_36963

   PIN FE_OFN71221_n_51388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.562 0.163 40.59 ;
      END
   END FE_OFN71221_n_51388

   PIN FE_OFN71870_n_49472
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.282 0.163 71.31 ;
      END
   END FE_OFN71870_n_49472

   PIN FE_OFN71874_n_48941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.602 0.163 63.63 ;
      END
   END FE_OFN71874_n_48941

   PIN FE_OFN71876_n_49492
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.442 0.163 67.47 ;
      END
   END FE_OFN71876_n_49492

   PIN FE_OFN71880_n_48888
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.098 76.637 2.126 76.8 ;
      END
   END FE_OFN71880_n_48888

   PIN FE_OFN71884_n_49381
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.098 76.637 2.126 76.8 ;
      END
   END FE_OFN71884_n_49381

   PIN FE_OFN71898_n_49468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.746 0.163 61.774 ;
      END
   END FE_OFN71898_n_49468

   PIN FE_OFN71900_n_48857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.834 0.163 54.862 ;
      END
   END FE_OFN71900_n_48857

   PIN FE_OFN71903_n_48879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.81 0.163 61.838 ;
      END
   END FE_OFN71903_n_48879

   PIN FE_OFN71950_n_49434
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.474 0.163 55.502 ;
      END
   END FE_OFN71950_n_49434

   PIN FE_OFN72307_n_35478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.546 0.163 34.574 ;
      END
   END FE_OFN72307_n_35478

   PIN FE_OFN72308_n_35478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.898 0.163 22.926 ;
      END
   END FE_OFN72308_n_35478

   PIN FE_OFN72343_n_40157
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.626 0.163 40.654 ;
      END
   END FE_OFN72343_n_40157

   PIN FE_OFN72353_n_34646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.522 0.163 17.55 ;
      END
   END FE_OFN72353_n_34646

   PIN FE_OFN72354_n_34646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 21.17 0.163 21.198 ;
      END
   END FE_OFN72354_n_34646

   PIN FE_OFN73017_n_35230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.346 0.163 31.374 ;
      END
   END FE_OFN73017_n_35230

   PIN FE_OFN74845_n_34783
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.962 0.163 14.99 ;
      END
   END FE_OFN74845_n_34783

   PIN FE_OFN74988_n_34728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.21 0.0 44.238 0.163 ;
      END
   END FE_OFN74988_n_34728

   PIN FE_OFN75036_n_39918
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 60.338 53.376 60.366 ;
      END
   END FE_OFN75036_n_39918

   PIN FE_OFN83546_n_36628
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.578 0.163 54.606 ;
      END
   END FE_OFN83546_n_36628

   PIN FE_OFN83569_n_36967
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.202 76.637 9.23 76.8 ;
      END
   END FE_OFN83569_n_36967

   PIN FE_OFN83591_n_36801
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 23.026 0.163 23.054 ;
      END
   END FE_OFN83591_n_36801

   PIN FE_OFN84427_n_48865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.922 0.163 31.95 ;
      END
   END FE_OFN84427_n_48865

   PIN FE_OFN84447_eq_15948_66_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.754 0.0 48.782 0.163 ;
      END
   END FE_OFN84447_eq_15948_66_n_18

   PIN FE_OFN84485_n_45279
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.386 0.163 46.414 ;
      END
   END FE_OFN84485_n_45279

   PIN FE_OFN84520_n_51062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.314 76.637 3.342 76.8 ;
      END
   END FE_OFN84520_n_51062

   PIN FE_OFN84522_n_51648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.258 76.637 6.286 76.8 ;
      END
   END FE_OFN84522_n_51648

   PIN FE_OFN84525_n_51588
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.034 76.637 2.062 76.8 ;
      END
   END FE_OFN84525_n_51588

   PIN FE_OFN84528_n_48932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.146 76.637 4.174 76.8 ;
      END
   END FE_OFN84528_n_48932

   PIN FE_OFN84547_n_51122
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.93 76.637 2.958 76.8 ;
      END
   END FE_OFN84547_n_51122

   PIN FE_OFN84549_n_51605
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.61 0.163 58.638 ;
      END
   END FE_OFN84549_n_51605

   PIN FE_OFN84711_n_48951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.402 0.163 60.43 ;
      END
   END FE_OFN84711_n_48951

   PIN FE_OFN84743_n_61607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 53.49 53.376 53.518 ;
      END
   END FE_OFN84743_n_61607

   PIN FE_OFN86863_n_34728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.45 0.163 14.478 ;
      END
   END FE_OFN86863_n_34728

   PIN FE_OFN87003_n_36103
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 57.842 53.376 57.87 ;
      END
   END FE_OFN87003_n_36103

   PIN FE_OFN97682_n_36483
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 52.082 53.376 52.11 ;
      END
   END FE_OFN97682_n_36483

   PIN FE_OFN97790_n_7079
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.426 76.637 29.454 76.8 ;
      END
   END FE_OFN97790_n_7079

   PIN FE_OFN98056_n_43238
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.586 0.163 57.614 ;
      END
   END FE_OFN98056_n_43238

   PIN FE_OFN98707_n_35230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.962 0.163 30.99 ;
      END
   END FE_OFN98707_n_35230

   PIN FE_RN_1121_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.826 0.163 51.854 ;
      END
   END FE_RN_1121_0

   PIN FE_RN_1136_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.418 0.0 26.446 0.163 ;
      END
   END FE_RN_1136_0

   PIN FE_RN_1694_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.914 0.163 28.942 ;
      END
   END FE_RN_1694_0

   PIN add_85566_69_n_36
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 61.17 53.376 61.198 ;
      END
   END add_85566_69_n_36

   PIN eq_15818_44_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.65 0.163 41.678 ;
      END
   END eq_15818_44_n_18

   PIN eq_15822_44_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.986 0.163 32.014 ;
      END
   END eq_15822_44_n_18

   PIN eq_15848_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.626 0.163 8.654 ;
      END
   END eq_15848_46_n_18

   PIN eq_15858_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.674 0.163 42.702 ;
      END
   END eq_15858_46_n_18

   PIN eq_15862_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 43.634 0.163 43.662 ;
      END
   END eq_15862_46_n_18

   PIN eq_15866_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.69 0.0 32.718 0.163 ;
      END
   END eq_15866_46_n_18

   PIN g2_m_5__3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.874 0.163 61.902 ;
      END
   END g2_m_5__3_

   PIN memread_edit_dist_g2_ln254_unr6_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.826 76.637 27.854 76.8 ;
      END
   END memread_edit_dist_g2_ln254_unr6_q_0_

   PIN memread_edit_dist_g2_ln254_unr6_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.938 76.637 45.966 76.8 ;
      END
   END memread_edit_dist_g2_ln254_unr6_q_3_

   PIN mux_g_ln477_q_117_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 47.282 53.376 47.31 ;
      END
   END mux_g_ln477_q_117_

   PIN mux_g_ln477_q_128_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 40.242 53.376 40.27 ;
      END
   END mux_g_ln477_q_128_

   PIN n_10566
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.354 76.637 18.382 76.8 ;
      END
   END n_10566

   PIN n_11993
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.162 0.163 58.19 ;
      END
   END n_11993

   PIN n_11994
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.034 0.163 66.062 ;
      END
   END n_11994

   PIN n_11995
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 65.522 53.376 65.55 ;
      END
   END n_11995

   PIN n_11997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.282 0.163 63.31 ;
      END
   END n_11997

   PIN n_11998
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.082 0.163 68.11 ;
      END
   END n_11998

   PIN n_11999
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 66.418 53.376 66.446 ;
      END
   END n_11999

   PIN n_12000
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.314 0.163 75.342 ;
      END
   END n_12000

   PIN n_12001
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 62.322 53.376 62.35 ;
      END
   END n_12001

   PIN n_12002
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.098 0.163 66.126 ;
      END
   END n_12002

   PIN n_12003
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 71.73 53.376 71.758 ;
      END
   END n_12003

   PIN n_12004
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.418 0.163 66.446 ;
      END
   END n_12004

   PIN n_12005
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 53.213 66.354 53.376 66.382 ;
      END
   END n_12005

   PIN n_12006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.986 0.163 72.014 ;
      END
   END n_12006

   PIN n_12026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.162 0.163 66.19 ;
      END
   END n_12026

   PIN n_12027
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.85 0.163 60.878 ;
      END
   END n_12027

   PIN n_12345
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 63.282 53.376 63.31 ;
      END
   END n_12345

   PIN n_12353
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.29 0.163 66.318 ;
      END
   END n_12353

   PIN n_12926
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.698 0.163 75.726 ;
      END
   END n_12926

   PIN n_12932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.762 0.163 75.79 ;
      END
   END n_12932

   PIN n_14365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 61.426 53.376 61.454 ;
      END
   END n_14365

   PIN n_14987
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.826 0.163 75.854 ;
      END
   END n_14987

   PIN n_15857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 68.722 53.376 68.75 ;
      END
   END n_15857

   PIN n_15877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 69.106 53.376 69.134 ;
      END
   END n_15877

   PIN n_17531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 66.034 53.376 66.062 ;
      END
   END n_17531

   PIN n_17902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 64.754 53.376 64.782 ;
      END
   END n_17902

   PIN n_18259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 63.09 53.376 63.118 ;
      END
   END n_18259

   PIN n_18380
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 66.162 53.376 66.19 ;
      END
   END n_18380

   PIN n_18657
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.466 0.082 68.494 ;
      END
   END n_18657

   PIN n_18826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.242 0.0 8.27 0.163 ;
      END
   END n_18826

   PIN n_21936
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 61.298 53.376 61.326 ;
      END
   END n_21936

   PIN n_2287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.346 0.163 71.374 ;
      END
   END n_2287

   PIN n_25366
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.474 0.163 31.502 ;
      END
   END n_25366

   PIN n_25372
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.842 0.163 25.87 ;
      END
   END n_25372

   PIN n_31455
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 57.906 53.376 57.934 ;
      END
   END n_31455

   PIN n_3429
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.642 76.637 46.67 76.8 ;
      END
   END n_3429

   PIN n_34414
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 43.506 0.163 43.534 ;
      END
   END n_34414

   PIN n_34611
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.154 0.082 15.182 ;
      END
   END n_34611

   PIN n_34613
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.642 0.082 22.67 ;
      END
   END n_34613

   PIN n_34614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.322 0.082 14.35 ;
      END
   END n_34614

   PIN n_34647
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.29 0.082 18.318 ;
      END
   END n_34647

   PIN n_34648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.738 0.082 34.766 ;
      END
   END n_34648

   PIN n_34649
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.978 0.163 29.006 ;
      END
   END n_34649

   PIN n_34684
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.842 0.163 33.87 ;
      END
   END n_34684

   PIN n_35083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 37.298 0.163 37.326 ;
      END
   END n_35083

   PIN n_35219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.346 0.163 39.374 ;
      END
   END n_35219

   PIN n_35229
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.242 0.082 32.27 ;
      END
   END n_35229

   PIN n_35231
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.33 0.082 25.358 ;
      END
   END n_35231

   PIN n_35232
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.69 0.082 8.718 ;
      END
   END n_35232

   PIN n_35448
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 30.258 0.163 30.286 ;
      END
   END n_35448

   PIN n_35471
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.13 0.082 14.158 ;
      END
   END n_35471

   PIN n_35472
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.834 0.163 22.862 ;
      END
   END n_35472

   PIN n_35475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 5.426 0.163 5.454 ;
      END
   END n_35475

   PIN n_35476
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.602 0.163 31.63 ;
      END
   END n_35476

   PIN n_35477
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.106 0.082 37.134 ;
      END
   END n_35477

   PIN n_35479
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.274 0.163 20.302 ;
      END
   END n_35479

   PIN n_35507
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.738 0.163 18.766 ;
      END
   END n_35507

   PIN n_35515
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.162 0.163 2.19 ;
      END
   END n_35515

   PIN n_35563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 23.41 0.082 23.438 ;
      END
   END n_35563

   PIN n_35567
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.354 0.082 18.382 ;
      END
   END n_35567

   PIN n_35590
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.042 0.163 29.07 ;
      END
   END n_35590

   PIN n_35722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.922 0.163 15.95 ;
      END
   END n_35722

   PIN n_35728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.89 0.163 11.918 ;
      END
   END n_35728

   PIN n_35774
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 18.93 53.376 18.958 ;
      END
   END n_35774

   PIN n_35775
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.65 0.163 25.678 ;
      END
   END n_35775

   PIN n_3604
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.322 76.637 14.35 76.8 ;
      END
   END n_3604

   PIN n_3608
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.418 76.637 18.446 76.8 ;
      END
   END n_3608

   PIN n_36089
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 60.402 53.376 60.43 ;
      END
   END n_36089

   PIN n_3612
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 70.386 0.163 70.414 ;
      END
   END n_3612

   PIN n_36199
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.794 53.376 31.822 ;
      END
   END n_36199

   PIN n_36776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 46.642 0.0 46.67 0.163 ;
      END
   END n_36776

   PIN n_36959
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.266 76.637 9.294 76.8 ;
      END
   END n_36959

   PIN n_37013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.178 76.637 32.206 76.8 ;
      END
   END n_37013

   PIN n_37017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 75.122 0.163 75.15 ;
      END
   END n_37017

   PIN n_37026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 54.002 53.376 54.03 ;
      END
   END n_37026

   PIN n_37033
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 57.714 53.376 57.742 ;
      END
   END n_37033

   PIN n_39567
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.186 0.163 43.214 ;
      END
   END n_39567

   PIN n_39579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 41.202 0.163 41.23 ;
      END
   END n_39579

   PIN n_39580
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.37 0.163 40.398 ;
      END
   END n_39580

   PIN n_39675
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.538 0.163 15.566 ;
      END
   END n_39675

   PIN n_39833
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.586 0.163 25.614 ;
      END
   END n_39833

   PIN n_39839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.466 0.163 28.494 ;
      END
   END n_39839

   PIN n_39854
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 18.226 53.376 18.254 ;
      END
   END n_39854

   PIN n_39882
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.154 0.163 63.182 ;
      END
   END n_39882

   PIN n_39911
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 50.802 53.376 50.83 ;
      END
   END n_39911

   PIN n_39920
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 34.61 53.376 34.638 ;
      END
   END n_39920

   PIN n_39965
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.01 0.163 33.038 ;
      END
   END n_39965

   PIN n_40114
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.058 0.163 35.086 ;
      END
   END n_40114

   PIN n_41399
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.09 0.163 23.118 ;
      END
   END n_41399

   PIN n_41410
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.322 0.163 38.35 ;
      END
   END n_41410

   PIN n_41424
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.994 0.163 43.022 ;
      END
   END n_41424

   PIN n_42305
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.674 0.163 18.702 ;
      END
   END n_42305

   PIN n_42524
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.178 0.0 32.206 0.163 ;
      END
   END n_42524

   PIN n_42707
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 1.97 53.376 1.998 ;
      END
   END n_42707

   PIN n_42987
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.002 0.163 38.03 ;
      END
   END n_42987

   PIN n_43058
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.666 0.163 31.694 ;
      END
   END n_43058

   PIN n_43098
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.73 0.163 31.758 ;
      END
   END n_43098

   PIN n_43116
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.538 0.163 31.566 ;
      END
   END n_43116

   PIN n_43142
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.202 0.163 41.23 ;
      END
   END n_43142

   PIN n_43174
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.058 0.163 3.086 ;
      END
   END n_43174

   PIN n_45172
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.946 0.163 8.974 ;
      END
   END n_45172

   PIN n_45277
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.386 0.163 38.414 ;
      END
   END n_45277

   PIN n_45524
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 28.594 0.163 28.622 ;
      END
   END n_45524

   PIN n_45825
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 5.938 53.376 5.966 ;
      END
   END n_45825

   PIN n_45972
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.61 0.163 18.638 ;
      END
   END n_45972

   PIN n_46005
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.714 0.163 25.742 ;
      END
   END n_46005

   PIN n_46166
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.378 0.163 11.406 ;
      END
   END n_46166

   PIN n_46167
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.442 0.163 11.47 ;
      END
   END n_46167

   PIN n_46192
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.474 0.0 23.502 0.163 ;
      END
   END n_46192

   PIN n_46540
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 29.042 53.376 29.07 ;
      END
   END n_46540

   PIN n_46555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 6.002 53.376 6.03 ;
      END
   END n_46555

   PIN n_46557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.842 0.0 17.87 0.163 ;
      END
   END n_46557

   PIN n_48369
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.65 0.163 57.678 ;
      END
   END n_48369

   PIN n_48630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 43.57 0.163 43.598 ;
      END
   END n_48630

   PIN n_48760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.242 0.0 32.27 0.163 ;
      END
   END n_48760

   PIN n_48784
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 6.066 53.376 6.094 ;
      END
   END n_48784

   PIN n_48790
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 14.45 53.376 14.478 ;
      END
   END n_48790

   PIN n_48801
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 14.514 53.376 14.542 ;
      END
   END n_48801

   PIN n_48882
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.738 0.0 18.766 0.163 ;
      END
   END n_48882

   PIN n_48894
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 46.194 0.163 46.222 ;
      END
   END n_48894

   PIN n_48907
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.242 0.163 72.27 ;
      END
   END n_48907

   PIN n_48913
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.89 0.163 51.918 ;
      END
   END n_48913

   PIN n_48927
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 52.53 0.163 52.558 ;
      END
   END n_48927

   PIN n_49353
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.218 0.163 15.246 ;
      END
   END n_49353

   PIN n_49364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.434 0.163 48.462 ;
      END
   END n_49364

   PIN n_49837
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 66.29 0.163 66.318 ;
      END
   END n_49837

   PIN n_5042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 32.242 0.163 32.27 ;
      END
   END n_5042

   PIN n_51039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.338 0.163 60.366 ;
      END
   END n_51039

   PIN n_51043
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 54.898 0.163 54.926 ;
      END
   END n_51043

   PIN n_51046
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.034 76.637 18.062 76.8 ;
      END
   END n_51046

   PIN n_51219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.77 0.163 54.798 ;
      END
   END n_51219

   PIN n_51577
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.538 0.163 63.566 ;
      END
   END n_51577

   PIN n_51584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.306 0.163 72.334 ;
      END
   END n_51584

   PIN n_51600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.346 0.163 63.374 ;
      END
   END n_51600

   PIN n_51640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.074 76.637 33.102 76.8 ;
      END
   END n_51640

   PIN n_51655
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.058 0.163 75.086 ;
      END
   END n_51655

   PIN n_51678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.098 0.163 2.126 ;
      END
   END n_51678

   PIN n_51711
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.466 0.163 60.494 ;
      END
   END n_51711

   PIN n_5226968_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 38.002 53.376 38.03 ;
      END
   END n_5226968_bar

   PIN n_58231
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 36.85 53.376 36.878 ;
      END
   END n_58231

   PIN n_58248
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 37.426 53.376 37.454 ;
      END
   END n_58248

   PIN n_58255
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 38.13 53.376 38.158 ;
      END
   END n_58255

   PIN n_58274
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 11.698 53.376 11.726 ;
      END
   END n_58274

   PIN n_58468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.858 53.376 31.886 ;
      END
   END n_58468

   PIN n_58771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 38.642 53.376 38.67 ;
      END
   END n_58771

   PIN n_60940
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.29 0.163 34.318 ;
      END
   END n_60940

   PIN n_61
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.018 76.637 12.046 76.8 ;
      END
   END n_61

   PIN n_61009
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.874 0.163 45.902 ;
      END
   END n_61009

   PIN n_61819
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.794 0.163 31.822 ;
      END
   END n_61819

   PIN n_65255
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.954 0.163 11.982 ;
      END
   END n_65255

   PIN n_65263
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.074 0.0 33.102 0.163 ;
      END
   END n_65263

   PIN n_65290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.114 76.637 32.142 76.8 ;
      END
   END n_65290

   PIN n_65302
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.058 76.637 35.086 76.8 ;
      END
   END n_65302

   PIN n_8376
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.818 0.163 64.846 ;
      END
   END n_8376

   PIN n_9348
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 66.226 53.376 66.254 ;
      END
   END n_9348

   PIN n_9349
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 69.17 53.376 69.198 ;
      END
   END n_9349

   PIN n_9350
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 68.082 53.376 68.11 ;
      END
   END n_9350

   PIN n_9351
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 68.146 53.376 68.174 ;
      END
   END n_9351

   PIN n_9353
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 68.402 53.376 68.43 ;
      END
   END n_9353

   PIN sub_14960_49_n_107
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.386 0.163 14.414 ;
      END
   END sub_14960_49_n_107

   PIN sub_14970_49_n_107
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.906 0.163 25.934 ;
      END
   END sub_14970_49_n_107

   PIN sub_14999_49_n_108
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 37.362 0.163 37.39 ;
      END
   END sub_14999_49_n_108

   PIN sub_15894_74_n_2572416
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.506 0.163 35.534 ;
      END
   END sub_15894_74_n_2572416

   PIN sub_ln263_unr104_z_3__4326697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.738 0.163 34.766 ;
      END
   END sub_ln263_unr104_z_3__4326697

   PIN sub_ln263_unr36_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.45 0.163 38.478 ;
      END
   END sub_ln263_unr36_z_6_

   PIN sub_ln263_unr52_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.722 0.163 36.75 ;
      END
   END sub_ln263_unr52_z_6_

   PIN ternarymux_ln49_0_unr7_z_0__4472252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 54.322 53.376 54.35 ;
      END
   END ternarymux_ln49_0_unr7_z_0__4472252

   PIN ternarymux_ln49_0_unr7_z_1__4472242
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 51.89 53.376 51.918 ;
      END
   END ternarymux_ln49_0_unr7_z_1__4472242

   PIN ternarymux_ln49_0_unr7_z_2__4472244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 54.962 53.376 54.99 ;
      END
   END ternarymux_ln49_0_unr7_z_2__4472244

   PIN FE_OCPN57641_sub_14990_49_n_2572016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.746 0.163 29.774 ;
      END
   END FE_OCPN57641_sub_14990_49_n_2572016

   PIN FE_OCPN57647_FE_OFN47241_n_6273_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.61 0.163 42.638 ;
      END
   END FE_OCPN57647_FE_OFN47241_n_6273_bar

   PIN FE_OCPN57979_FE_OFN47238_mux_k_ln251_z_5__4323813_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.714 0.163 41.742 ;
      END
   END FE_OCPN57979_FE_OFN47238_mux_k_ln251_z_5__4323813_bar

   PIN FE_OCPN58925_n_35465
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.106 0.163 45.134 ;
      END
   END FE_OCPN58925_n_35465

   PIN FE_OCPN59173_add_15054_37_n_30
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.842 0.163 25.87 ;
      END
   END FE_OCPN59173_add_15054_37_n_30

   PIN FE_OCPN61716_n_25369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.482 0.163 34.51 ;
      END
   END FE_OCPN61716_n_25369

   PIN FE_OCPN62290_FE_OFN54291_sub_15040_54_n_2572501
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.586 0.163 25.614 ;
      END
   END FE_OCPN62290_FE_OFN54291_sub_15040_54_n_2572501

   PIN FE_OCPN62338_n_65283
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 28.85 53.376 28.878 ;
      END
   END FE_OCPN62338_n_65283

   PIN FE_OCPN63182_n_34649
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.594 0.082 28.622 ;
      END
   END FE_OCPN63182_n_34649

   PIN FE_OCPN63193_n_35226
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 36.722 0.163 36.75 ;
      END
   END FE_OCPN63193_n_35226

   PIN FE_OCPN63292_sub_15039_54_n_48
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.106 0.163 29.134 ;
      END
   END FE_OCPN63292_sub_15039_54_n_48

   PIN FE_OCPN63324_n_35588
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.482 0.163 26.51 ;
      END
   END FE_OCPN63324_n_35588

   PIN FE_OCPN63391_FE_OFN37146_sub_15016_49_n_98_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.146 0.163 20.174 ;
      END
   END FE_OCPN63391_FE_OFN37146_sub_15016_49_n_98_bar

   PIN FE_OCPN63717_FE_OFN38588_mux_k_ln251_z_6__4323808_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.434 0.163 40.462 ;
      END
   END FE_OCPN63717_FE_OFN38588_mux_k_ln251_z_6__4323808_bar

   PIN FE_OCPN63732_n_34650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.066 0.163 22.094 ;
      END
   END FE_OCPN63732_n_34650

   PIN FE_OCPN63734_n_34650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.794 0.082 15.822 ;
      END
   END FE_OCPN63734_n_34650

   PIN FE_OCPN63741_n_34677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.402 0.163 28.43 ;
      END
   END FE_OCPN63741_n_34677

   PIN FE_OCPN99275_n_31308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.522 76.637 49.55 76.8 ;
      END
   END FE_OCPN99275_n_31308

   PIN FE_OCP_RBN77513_n_58100
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 8.69 53.376 8.718 ;
      END
   END FE_OCP_RBN77513_n_58100

   PIN FE_OFN27525_n_36175
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.41 0.163 63.438 ;
      END
   END FE_OFN27525_n_36175

   PIN FE_OFN27527_n_36461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.938 76.637 37.966 76.8 ;
      END
   END FE_OFN27527_n_36461

   PIN FE_OFN27529_n_36817
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.65 0.163 57.678 ;
      END
   END FE_OFN27529_n_36817

   PIN FE_OFN27719_n_36831
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 43.122 53.376 43.15 ;
      END
   END FE_OFN27719_n_36831

   PIN FE_OFN27721_n_36822
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 37.042 53.376 37.07 ;
      END
   END FE_OFN27721_n_36822

   PIN FE_OFN27723_n_36770
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 41.97 53.376 41.998 ;
      END
   END FE_OFN27723_n_36770

   PIN FE_OFN27736_n_36719
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 66.354 53.376 66.382 ;
      END
   END FE_OFN27736_n_36719

   PIN FE_OFN27941_n_36634
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.594 76.637 44.622 76.8 ;
      END
   END FE_OFN27941_n_36634

   PIN FE_OFN27988_n_36594
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.762 76.637 43.79 76.8 ;
      END
   END FE_OFN27988_n_36594

   PIN FE_OFN28005_n_36578
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.482 76.637 26.51 76.8 ;
      END
   END FE_OFN28005_n_36578

   PIN FE_OFN28007_n_36087
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.962 76.637 14.99 76.8 ;
      END
   END FE_OFN28007_n_36087

   PIN FE_OFN28009_n_36576
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.898 76.637 14.926 76.8 ;
      END
   END FE_OFN28009_n_36576

   PIN FE_OFN28011_n_36573
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.498 76.637 24.526 76.8 ;
      END
   END FE_OFN28011_n_36573

   PIN FE_OFN28149_n_36991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.162 76.637 2.19 76.8 ;
      END
   END FE_OFN28149_n_36991

   PIN FE_OFN28263_n_36480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.322 76.637 6.35 76.8 ;
      END
   END FE_OFN28263_n_36480

   PIN FE_OFN28266_n_37062
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 49.01 0.163 49.038 ;
      END
   END FE_OFN28266_n_37062

   PIN FE_OFN28302_n_36267
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.586 76.637 49.614 76.8 ;
      END
   END FE_OFN28302_n_36267

   PIN FE_OFN29813_n_59339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.73 76.718 31.758 76.8 ;
      END
   END FE_OFN29813_n_59339

   PIN FE_OFN30059_n_34783
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 34.546 53.376 34.574 ;
      END
   END FE_OFN30059_n_34783

   PIN FE_OFN30063_n_39931
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.714 0.163 57.742 ;
      END
   END FE_OFN30063_n_39931

   PIN FE_OFN30374_n_34771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 46.642 76.718 46.67 76.8 ;
      END
   END FE_OFN30374_n_34771

   PIN FE_OFN30391_n_34771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 47.09 53.376 47.118 ;
      END
   END FE_OFN30391_n_34771

   PIN FE_OFN30393_n_34771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.738 76.718 34.766 76.8 ;
      END
   END FE_OFN30393_n_34771

   PIN FE_OFN30500_n_34778
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 40.946 53.376 40.974 ;
      END
   END FE_OFN30500_n_34778

   PIN FE_OFN30777_n_34754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.746 76.718 37.774 76.8 ;
      END
   END FE_OFN30777_n_34754

   PIN FE_OFN33694_n_871
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.722 76.637 20.75 76.8 ;
      END
   END FE_OFN33694_n_871

   PIN FE_OFN33863_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.506 0.163 75.534 ;
      END
   END FE_OFN33863_n_71

   PIN FE_OFN33942_n_93
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.322 76.637 6.35 76.8 ;
      END
   END FE_OFN33942_n_93

   PIN FE_OFN34078_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.202 76.637 9.23 76.8 ;
      END
   END FE_OFN34078_n_87

   PIN FE_OFN34099_n_86
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.882 76.637 24.91 76.8 ;
      END
   END FE_OFN34099_n_86

   PIN FE_OFN34189_n_82
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.402 0.163 44.43 ;
      END
   END FE_OFN34189_n_82

   PIN FE_OFN34490_n_224
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.802 0.163 50.83 ;
      END
   END FE_OFN34490_n_224

   PIN FE_OFN34615_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 40.562 53.376 40.59 ;
      END
   END FE_OFN34615_n_223

   PIN FE_OFN35134_n_61599
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.642 0.163 54.67 ;
      END
   END FE_OFN35134_n_61599

   PIN FE_OFN35392_n_43250
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.362 0.163 37.39 ;
      END
   END FE_OFN35392_n_43250

   PIN FE_OFN35421_eq_15766_42_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.786 0.0 20.814 0.163 ;
      END
   END FE_OFN35421_eq_15766_42_n_18

   PIN FE_OFN35722_n_49478
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.09 0.0 7.118 0.163 ;
      END
   END FE_OFN35722_n_49478

   PIN FE_OFN35745_n_60966
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.466 0.0 12.494 0.163 ;
      END
   END FE_OFN35745_n_60966

   PIN FE_OFN36439_n_43089
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.122 0.163 3.15 ;
      END
   END FE_OFN36439_n_43089

   PIN FE_OFN36449_n_39997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.738 0.163 18.766 ;
      END
   END FE_OFN36449_n_39997

   PIN FE_OFN36464_n_43125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.346 0.0 23.374 0.163 ;
      END
   END FE_OFN36464_n_43125

   PIN FE_OFN36476_n_39651
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.426 0.163 5.454 ;
      END
   END FE_OFN36476_n_39651

   PIN FE_OFN36503_n_48575
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 5.362 53.376 5.39 ;
      END
   END FE_OFN36503_n_48575

   PIN FE_OFN36505_n_43150
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.41 0.0 15.438 0.163 ;
      END
   END FE_OFN36505_n_43150

   PIN FE_OFN36515_n_45481
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.722 0.163 4.75 ;
      END
   END FE_OFN36515_n_45481

   PIN FE_OFN36569_n_34614
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END FE_OFN36569_n_34614

   PIN FE_OFN36584_n_51062
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.57 0.0 3.598 0.163 ;
      END
   END FE_OFN36584_n_51062

   PIN FE_OFN36712_n_35722
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.602 0.163 15.63 ;
      END
   END FE_OFN36712_n_35722

   PIN FE_OFN36738_n_45529
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.906 0.163 1.934 ;
      END
   END FE_OFN36738_n_45529

   PIN FE_OFN36754_n_35564
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 23.282 0.163 23.31 ;
      END
   END FE_OFN36754_n_35564

   PIN FE_OFN36782_n_43330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.202 0.0 9.23 0.163 ;
      END
   END FE_OFN36782_n_43330

   PIN FE_OFN36821_n_48932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.506 0.0 3.534 0.163 ;
      END
   END FE_OFN36821_n_48932

   PIN FE_OFN37107_n_39853
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 6.13 53.376 6.158 ;
      END
   END FE_OFN37107_n_39853

   PIN FE_OFN37260_n_45839
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.562 0.163 8.59 ;
      END
   END FE_OFN37260_n_45839

   PIN FE_OFN37689_n_45290
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.242 0.0 32.27 0.163 ;
      END
   END FE_OFN37689_n_45290

   PIN FE_OFN37713_n_45400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.922 0.0 23.95 0.163 ;
      END
   END FE_OFN37713_n_45400

   PIN FE_OFN37718_n_39688
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.762 0.163 11.79 ;
      END
   END FE_OFN37718_n_39688

   PIN FE_OFN38279_sub_15035_54_n_74
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.65 0.163 25.678 ;
      END
   END FE_OFN38279_sub_15035_54_n_74

   PIN FE_OFN38497_n_42702
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.162 0.163 18.19 ;
      END
   END FE_OFN38497_n_42702

   PIN FE_OFN40808_n_35230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 30.13 0.082 30.158 ;
      END
   END FE_OFN40808_n_35230

   PIN FE_OFN40809_n_35230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.17 0.163 29.198 ;
      END
   END FE_OFN40809_n_35230

   PIN FE_OFN41487_sub_15027_54_n_55
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.522 0.163 41.55 ;
      END
   END FE_OFN41487_sub_15027_54_n_55

   PIN FE_OFN41911_n_227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.442 0.163 75.47 ;
      END
   END FE_OFN41911_n_227

   PIN FE_OFN41974_n_228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.538 0.163 47.566 ;
      END
   END FE_OFN41974_n_228

   PIN FE_OFN41984_n_228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 48.818 53.376 48.846 ;
      END
   END FE_OFN41984_n_228

   PIN FE_OFN42379_n_44
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.722 76.637 20.75 76.8 ;
      END
   END FE_OFN42379_n_44

   PIN FE_OFN42673_n_16
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.762 76.637 43.79 76.8 ;
      END
   END FE_OFN42673_n_16

   PIN FE_OFN42800_n_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.05 76.637 32.078 76.8 ;
      END
   END FE_OFN42800_n_11

   PIN FE_OFN42823_n_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.554 76.637 37.582 76.8 ;
      END
   END FE_OFN42823_n_10

   PIN FE_OFN43021_n_35315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 75.186 53.376 75.214 ;
      END
   END FE_OFN43021_n_35315

   PIN FE_OFN43045_n_35324
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 46.962 53.376 46.99 ;
      END
   END FE_OFN43045_n_35324

   PIN FE_OFN43227_n_35284
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.986 76.637 32.014 76.8 ;
      END
   END FE_OFN43227_n_35284

   PIN FE_OFN43246_n_35279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.058 76.637 35.086 76.8 ;
      END
   END FE_OFN43246_n_35279

   PIN FE_OFN43814_n_67218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.146 76.718 12.174 76.8 ;
      END
   END FE_OFN43814_n_67218

   PIN FE_OFN47463_sub_14941_55_n_80
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.778 0.163 25.806 ;
      END
   END FE_OFN47463_sub_14941_55_n_80

   PIN FE_OFN47468_sub_15027_54_n_55
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.986 0.163 40.014 ;
      END
   END FE_OFN47468_sub_15027_54_n_55

   PIN FE_OFN48046_sub_14960_49_n_142
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.826 0.163 11.854 ;
      END
   END FE_OFN48046_sub_14960_49_n_142

   PIN FE_OFN48509_n_59356
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 25.202 53.376 25.23 ;
      END
   END FE_OFN48509_n_59356

   PIN FE_OFN49847_n_77
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.402 76.637 28.43 76.8 ;
      END
   END FE_OFN49847_n_77

   PIN FE_OFN49963_n_48908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.786 0.163 68.814 ;
      END
   END FE_OFN49963_n_48908

   PIN FE_OFN50044_n_49472
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.474 0.163 63.502 ;
      END
   END FE_OFN50044_n_49472

   PIN FE_OFN50045_n_51588
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 5.874 0.163 5.902 ;
      END
   END FE_OFN50045_n_51588

   PIN FE_OFN50048_n_51648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.322 0.0 6.35 0.163 ;
      END
   END FE_OFN50048_n_51648

   PIN FE_OFN50217_n_51418
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.722 0.0 20.75 0.163 ;
      END
   END FE_OFN50217_n_51418

   PIN FE_OFN50653_n_58010
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 5.874 53.376 5.902 ;
      END
   END FE_OFN50653_n_58010

   PIN FE_OFN50871_n_35287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 48.242 53.376 48.27 ;
      END
   END FE_OFN50871_n_35287

   PIN FE_OFN54182_n_57313
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.362 0.0 45.39 0.163 ;
      END
   END FE_OFN54182_n_57313

   PIN FE_OFN54227_n_57317
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 8.626 53.376 8.654 ;
      END
   END FE_OFN54227_n_57317

   PIN FE_OFN54578_n_21110
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 47.474 53.376 47.502 ;
      END
   END FE_OFN54578_n_21110

   PIN FE_OFN64099_n_55937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.818 0.163 48.846 ;
      END
   END FE_OFN64099_n_55937

   PIN FE_OFN71220_n_51388
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.57 0.0 43.598 0.163 ;
      END
   END FE_OFN71220_n_51388

   PIN FE_OFN71873_n_48941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.714 0.163 57.742 ;
      END
   END FE_OFN71873_n_48941

   PIN FE_OFN71875_n_49492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.594 0.163 60.622 ;
      END
   END FE_OFN71875_n_49492

   PIN FE_OFN71879_n_48888
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.53 0.163 60.558 ;
      END
   END FE_OFN71879_n_48888

   PIN FE_OFN71883_n_49381
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.41 0.163 63.438 ;
      END
   END FE_OFN71883_n_49381

   PIN FE_OFN71949_n_49434
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.282 0.163 55.31 ;
      END
   END FE_OFN71949_n_49434

   PIN FE_OFN72112_n_45317
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 2.034 53.376 2.062 ;
      END
   END FE_OFN72112_n_45317

   PIN FE_OFN72158_n_43112
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.042 0.0 21.07 0.163 ;
      END
   END FE_OFN72158_n_43112

   PIN FE_OFN72170_n_42489
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 15.602 53.376 15.63 ;
      END
   END FE_OFN72170_n_42489

   PIN FE_OFN72809_sub_14939_54_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.058 0.163 19.086 ;
      END
   END FE_OFN72809_sub_14939_54_n_87

   PIN FE_OFN73560_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.602 76.637 39.63 76.8 ;
      END
   END FE_OFN73560_n_50

   PIN FE_OFN73816_n_234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.362 76.637 29.39 76.8 ;
      END
   END FE_OFN73816_n_234

   PIN FE_OFN74055_ternarymux_ln49_0_unr7_z_3__4472243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 63.218 53.376 63.246 ;
      END
   END FE_OFN74055_ternarymux_ln49_0_unr7_z_3__4472243

   PIN FE_OFN74157_n_883
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.706 0.163 54.734 ;
      END
   END FE_OFN74157_n_883

   PIN FE_OFN74165_n_876
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.698 0.0 11.726 0.163 ;
      END
   END FE_OFN74165_n_876

   PIN FE_OFN74186_n_875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.138 0.0 9.166 0.163 ;
      END
   END FE_OFN74186_n_875

   PIN FE_OFN74237_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.434 0.082 72.462 ;
      END
   END FE_OFN74237_n_223

   PIN FE_OFN74738_n_526
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.082 76.637 12.11 76.8 ;
      END
   END FE_OFN74738_n_526

   PIN FE_OFN74885_n_34782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.434 76.637 40.462 76.8 ;
      END
   END FE_OFN74885_n_34782

   PIN FE_OFN74896_n_34780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 43.826 53.376 43.854 ;
      END
   END FE_OFN74896_n_34780

   PIN FE_OFN74982_n_34728
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 54.898 53.376 54.926 ;
      END
   END FE_OFN74982_n_34728

   PIN FE_OFN75096_n_34784
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.138 76.637 9.166 76.8 ;
      END
   END FE_OFN75096_n_34784

   PIN FE_OFN75341_n_35324
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.242 76.637 32.27 76.8 ;
      END
   END FE_OFN75341_n_35324

   PIN FE_OFN75380_n_35283
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.298 76.637 29.326 76.8 ;
      END
   END FE_OFN75380_n_35283

   PIN FE_OFN75718_FE_OCPN56136_n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.562 0.163 40.59 ;
      END
   END FE_OFN75718_FE_OCPN56136_n_35331

   PIN FE_OFN75726_n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 71.346 0.163 71.374 ;
      END
   END FE_OFN75726_n_35331

   PIN FE_OFN79437_n_57254
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.882 0.0 40.91 0.163 ;
      END
   END FE_OFN79437_n_57254

   PIN FE_OFN83573_n_36956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 46.322 53.376 46.35 ;
      END
   END FE_OFN83573_n_36956

   PIN FE_OFN84709_n_43175
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.178 0.163 40.206 ;
      END
   END FE_OFN84709_n_43175

   PIN FE_OFN84938_n_7043
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.21 0.163 52.238 ;
      END
   END FE_OFN84938_n_7043

   PIN FE_OFN85149_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.538 76.637 23.566 76.8 ;
      END
   END FE_OFN85149_n_222

   PIN FE_OFN85189_n_226
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 36.018 53.376 36.046 ;
      END
   END FE_OFN85189_n_226

   PIN FE_OFN86333_n_4990
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 71.922 0.163 71.95 ;
      END
   END FE_OFN86333_n_4990

   PIN FE_OFN86459_n_7776
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 74.994 0.163 75.022 ;
      END
   END FE_OFN86459_n_7776

   PIN FE_OFN86874_n_34728
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 54.578 53.376 54.606 ;
      END
   END FE_OFN86874_n_34728

   PIN FE_OFN86916_n_34778
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 48.37 53.376 48.398 ;
      END
   END FE_OFN86916_n_34778

   PIN FE_OFN87971_n_35278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.938 76.637 37.966 76.8 ;
      END
   END FE_OFN87971_n_35278

   PIN FE_OFN90264_n_57193
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 23.282 53.376 23.31 ;
      END
   END FE_OFN90264_n_57193

   PIN FE_OFN93509_n_57220
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 34.162 53.376 34.19 ;
      END
   END FE_OFN93509_n_57220

   PIN FE_OFN95954_n_57193
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 26.034 53.376 26.062 ;
      END
   END FE_OFN95954_n_57193

   PIN FE_OFN97666_n_36632
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.914 76.637 36.942 76.8 ;
      END
   END FE_OFN97666_n_36632

   PIN FE_OFN97681_n_36483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 54.834 0.163 54.862 ;
      END
   END FE_OFN97681_n_36483

   PIN FE_OFN98055_n_43238
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.418 0.163 34.446 ;
      END
   END FE_OFN98055_n_43238

   PIN FE_OFN98229_n_865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.698 0.163 51.726 ;
      END
   END FE_OFN98229_n_865

   PIN FE_RN_1119_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.066 0.163 46.094 ;
      END
   END FE_RN_1119_0

   PIN FE_RN_1120_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.522 0.163 49.55 ;
      END
   END FE_RN_1120_0

   PIN b_in_16_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 75.122 53.376 75.15 ;
      END
   END b_in_16_2

   PIN b_in_16_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 53.213 49.074 53.376 49.102 ;
      END
   END b_in_16_3

   PIN b_in_18_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 60.658 53.376 60.686 ;
      END
   END b_in_18_1

   PIN b_in_18_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.378 76.637 35.406 76.8 ;
      END
   END b_in_18_2

   PIN b_in_22_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 53.213 46.194 53.376 46.222 ;
      END
   END b_in_22_0

   PIN b_in_22_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 53.213 63.474 53.376 63.502 ;
      END
   END b_in_22_2

   PIN b_in_22_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 46.13 53.376 46.158 ;
      END
   END b_in_22_3

   PIN b_in_26_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 53.213 70.386 53.376 70.414 ;
      END
   END b_in_26_1

   PIN b_in_26_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 53.213 43.506 53.376 43.534 ;
      END
   END b_in_26_3

   PIN b_in_29_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 53.213 46.066 53.376 46.094 ;
      END
   END b_in_29_1

   PIN b_in_32_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 53.213 40.434 53.376 40.462 ;
      END
   END b_in_32_0

   PIN eq_15778_44_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 49.138 0.163 49.166 ;
      END
   END eq_15778_44_n_18

   PIN eq_15782_44_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.018 0.0 12.046 0.163 ;
      END
   END eq_15782_44_n_18

   PIN eq_15784_44_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 45.042 53.376 45.07 ;
      END
   END eq_15784_44_n_18

   PIN g2_q8_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 61.362 53.376 61.39 ;
      END
   END g2_q8_2_

   PIN g2_q8_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 66.29 53.376 66.318 ;
      END
   END g2_q8_3_

   PIN gt_16017_52_n_89
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.258 0.163 38.286 ;
      END
   END gt_16017_52_n_89

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.122 0.082 51.15 ;
      END
   END ispd_clk

   PIN memread_edit_dist_g2_ln254_unr7_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 57.65 53.376 57.678 ;
      END
   END memread_edit_dist_g2_ln254_unr7_q_4_

   PIN memread_edit_dist_g2_ln254_unr7_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 57.778 53.376 57.806 ;
      END
   END memread_edit_dist_g2_ln254_unr7_q_6_

   PIN memread_edit_dist_g2_ln254_unr7_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 57.586 53.376 57.614 ;
      END
   END memread_edit_dist_g2_ln254_unr7_q_7_

   PIN memread_edit_dist_g2_ln254_unr8_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 43.89 53.376 43.918 ;
      END
   END memread_edit_dist_g2_ln254_unr8_q_11_

   PIN memread_edit_dist_g2_ln254_unr8_q_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 34.674 53.376 34.702 ;
      END
   END memread_edit_dist_g2_ln254_unr8_q_9_

   PIN mux_g_ln477_q_65_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.274 0.163 68.302 ;
      END
   END mux_g_ln477_q_65_

   PIN mux_k_ln251_z_7__4323810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 22.834 0.163 22.862 ;
      END
   END mux_k_ln251_z_7__4323810

   PIN n_11915
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.186 0.082 75.214 ;
      END
   END n_11915

   PIN n_12782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 63.154 53.376 63.182 ;
      END
   END n_12782

   PIN n_14602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.378 0.163 75.406 ;
      END
   END n_14602

   PIN n_15146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 65.138 53.376 65.166 ;
      END
   END n_15146

   PIN n_15147
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 65.01 53.376 65.038 ;
      END
   END n_15147

   PIN n_18127
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 69.042 53.376 69.07 ;
      END
   END n_18127

   PIN n_18128
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 66.098 53.376 66.126 ;
      END
   END n_18128

   PIN n_18558
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.922 0.163 71.95 ;
      END
   END n_18558

   PIN n_18559
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.138 0.163 65.166 ;
      END
   END n_18559

   PIN n_18725
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.178 0.163 72.206 ;
      END
   END n_18725

   PIN n_18732
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.978 0.163 69.006 ;
      END
   END n_18732

   PIN n_18789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.218 0.163 63.246 ;
      END
   END n_18789

   PIN n_18799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.226 0.163 66.254 ;
      END
   END n_18799

   PIN n_18800
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.114 0.163 72.142 ;
      END
   END n_18800

   PIN n_18801
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.074 0.163 65.102 ;
      END
   END n_18801

   PIN n_18802
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.722 0.163 68.75 ;
      END
   END n_18802

   PIN n_18803
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.01 0.163 65.038 ;
      END
   END n_18803

   PIN n_18804
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.21 0.163 68.238 ;
      END
   END n_18804

   PIN n_18805
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.522 0.163 57.55 ;
      END
   END n_18805

   PIN n_2103
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 43.762 53.376 43.79 ;
      END
   END n_2103

   PIN n_21081
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.642 0.0 6.67 0.163 ;
      END
   END n_21081

   PIN n_21433
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 45.682 0.163 45.71 ;
      END
   END n_21433

   PIN n_22021
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 61.234 53.376 61.262 ;
      END
   END n_22021

   PIN n_25369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.682 0.163 29.71 ;
      END
   END n_25369

   PIN n_25529
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.322 0.163 14.35 ;
      END
   END n_25529

   PIN n_31306
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 54.77 53.376 54.798 ;
      END
   END n_31306

   PIN n_3207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 40.178 53.376 40.206 ;
      END
   END n_3207

   PIN n_34362
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.922 0.163 39.95 ;
      END
   END n_34362

   PIN n_34472
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.458 0.163 25.486 ;
      END
   END n_34472

   PIN n_34609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.018 0.163 20.046 ;
      END
   END n_34609

   PIN n_34612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 28.466 0.082 28.494 ;
      END
   END n_34612

   PIN n_34634
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.994 0.163 19.022 ;
      END
   END n_34634

   PIN n_34645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.05 0.163 40.078 ;
      END
   END n_34645

   PIN n_34646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 27.122 0.163 27.15 ;
      END
   END n_34646

   PIN n_35217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.282 0.163 39.31 ;
      END
   END n_35217

   PIN n_35218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.194 0.163 38.222 ;
      END
   END n_35218

   PIN n_35228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 17.202 0.163 17.23 ;
      END
   END n_35228

   PIN n_35247
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.818 0.082 8.846 ;
      END
   END n_35247

   PIN n_35259
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.546 0.163 34.574 ;
      END
   END n_35259

   PIN n_35458
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.61 0.163 34.638 ;
      END
   END n_35458

   PIN n_35468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.034 0.163 2.062 ;
      END
   END n_35468

   PIN n_35499
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.442 0.163 19.47 ;
      END
   END n_35499

   PIN n_35514
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.618 0.163 5.646 ;
      END
   END n_35514

   PIN n_35556
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.866 0.163 34.894 ;
      END
   END n_35556

   PIN n_35613
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.874 0.163 5.902 ;
      END
   END n_35613

   PIN n_35675
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.442 0.163 35.47 ;
      END
   END n_35675

   PIN n_3606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.634 0.163 51.662 ;
      END
   END n_3606

   PIN n_3607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.506 0.163 11.534 ;
      END
   END n_3607

   PIN n_3610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.298 0.0 21.326 0.163 ;
      END
   END n_3610

   PIN n_36155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.986 76.637 24.014 76.8 ;
      END
   END n_36155

   PIN n_36176
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.362 76.637 13.39 76.8 ;
      END
   END n_36176

   PIN n_36231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.002 76.637 14.03 76.8 ;
      END
   END n_36231

   PIN n_36631
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.634 76.637 35.662 76.8 ;
      END
   END n_36631

   PIN n_36739
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.698 76.637 43.726 76.8 ;
      END
   END n_36739

   PIN n_36801
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 33.522 53.376 33.55 ;
      END
   END n_36801

   PIN n_39564
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.93 0.163 18.958 ;
      END
   END n_39564

   PIN n_39617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.37 0.163 40.398 ;
      END
   END n_39617

   PIN n_39641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.362 0.163 5.39 ;
      END
   END n_39641

   PIN n_39644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.97 0.163 1.998 ;
      END
   END n_39644

   PIN n_39646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.546 0.163 26.574 ;
      END
   END n_39646

   PIN n_39648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.554 0.163 5.582 ;
      END
   END n_39648

   PIN n_39682
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.258 0.163 14.286 ;
      END
   END n_39682

   PIN n_39687
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.754 0.082 8.782 ;
      END
   END n_39687

   PIN n_39918
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.738 76.637 42.766 76.8 ;
      END
   END n_39918

   PIN n_40005
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.082 0.163 20.11 ;
      END
   END n_40005

   PIN n_40121
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.674 0.163 18.702 ;
      END
   END n_40121

   PIN n_40134
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.01 0.163 17.038 ;
      END
   END n_40134

   PIN n_40243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.722 0.163 28.75 ;
      END
   END n_40243

   PIN n_41327
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.962 0.163 14.99 ;
      END
   END n_41327

   PIN n_42466
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 22.898 0.163 22.926 ;
      END
   END n_42466

   PIN n_42535
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.962 0.163 22.99 ;
      END
   END n_42535

   PIN n_42576
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.754 0.163 48.782 ;
      END
   END n_42576

   PIN n_43051
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.53 0.163 12.558 ;
      END
   END n_43051

   PIN n_43053
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.762 0.0 27.79 0.163 ;
      END
   END n_43053

   PIN n_43108
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.01 0.163 49.038 ;
      END
   END n_43108

   PIN n_43183
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.114 0.163 40.142 ;
      END
   END n_43183

   PIN n_43245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.386 0.0 22.414 0.163 ;
      END
   END n_43245

   PIN n_43247
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.242 0.163 40.27 ;
      END
   END n_43247

   PIN n_43262
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.714 0.163 25.742 ;
      END
   END n_43262

   PIN n_45279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.746 0.163 45.774 ;
      END
   END n_45279

   PIN n_45298
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.538 0.0 23.566 0.163 ;
      END
   END n_45298

   PIN n_45350
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.562 0.163 8.59 ;
      END
   END n_45350

   PIN n_45382
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.682 0.163 45.71 ;
      END
   END n_45382

   PIN n_45483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 18.162 53.376 18.19 ;
      END
   END n_45483

   PIN n_45488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.162 0.163 18.19 ;
      END
   END n_45488

   PIN n_46118
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.658 0.0 20.686 0.163 ;
      END
   END n_46118

   PIN n_46120
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.946 0.163 48.974 ;
      END
   END n_46120

   PIN n_46121
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.962 0.163 46.99 ;
      END
   END n_46121

   PIN n_46176
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 37.618 0.163 37.646 ;
      END
   END n_46176

   PIN n_46186
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.466 0.163 44.494 ;
      END
   END n_46186

   PIN n_468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 53.298 53.376 53.326 ;
      END
   END n_468

   PIN n_48346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.546 0.163 42.574 ;
      END
   END n_48346

   PIN n_48398
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.778 0.163 41.806 ;
      END
   END n_48398

   PIN n_48568
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.882 0.163 48.91 ;
      END
   END n_48568

   PIN n_48648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.13 0.163 38.158 ;
      END
   END n_48648

   PIN n_48764
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 22.962 0.163 22.99 ;
      END
   END n_48764

   PIN n_48806
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.306 0.163 40.334 ;
      END
   END n_48806

   PIN n_48859
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.322 0.163 62.35 ;
      END
   END n_48859

   PIN n_48865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.074 0.163 17.102 ;
      END
   END n_48865

   PIN n_48868
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.146 0.163 52.174 ;
      END
   END n_48868

   PIN n_48879
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.122 0.163 43.15 ;
      END
   END n_48879

   PIN n_48902
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.306 0.163 48.334 ;
      END
   END n_48902

   PIN n_48951
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.354 0.163 34.382 ;
      END
   END n_48951

   PIN n_49060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.882 0.163 8.91 ;
      END
   END n_49060

   PIN n_49063
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.466 0.163 12.494 ;
      END
   END n_49063

   PIN n_49214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.058 0.163 43.086 ;
      END
   END n_49214

   PIN n_49324
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.226 0.163 34.254 ;
      END
   END n_49324

   PIN n_49413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.298 0.163 37.326 ;
      END
   END n_49413

   PIN n_49468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.722 0.163 52.75 ;
      END
   END n_49468

   PIN n_49480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.978 0.163 13.006 ;
      END
   END n_49480

   PIN n_4992
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.314 76.637 27.342 76.8 ;
      END
   END n_4992

   PIN n_4999
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.682 0.163 61.71 ;
      END
   END n_4999

   PIN n_51064
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.482 0.163 58.51 ;
      END
   END n_51064

   PIN n_51122
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.666 0.163 31.694 ;
      END
   END n_51122

   PIN n_51575
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.994 0.163 3.022 ;
      END
   END n_51575

   PIN n_51605
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.602 0.163 31.63 ;
      END
   END n_51605

   PIN n_5223120_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.242 0.163 48.27 ;
      END
   END n_5223120_bar

   PIN n_5226969_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.234 0.163 37.262 ;
      END
   END n_5226969_bar

   PIN n_55934
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.946 0.163 48.974 ;
      END
   END n_55934

   PIN n_55936
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.042 0.163 45.07 ;
      END
   END n_55936

   PIN n_56252
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 46.13 0.163 46.158 ;
      END
   END n_56252

   PIN n_57047
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.754 0.0 24.782 0.163 ;
      END
   END n_57047

   PIN n_57053
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 12.146 0.163 12.174 ;
      END
   END n_57053

   PIN n_57311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 11.762 53.376 11.79 ;
      END
   END n_57311

   PIN n_57315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 8.562 53.376 8.59 ;
      END
   END n_57315

   PIN n_57327
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 8.754 53.376 8.782 ;
      END
   END n_57327

   PIN n_57353
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.482 0.0 26.51 0.163 ;
      END
   END n_57353

   PIN n_57645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.962 0.0 14.99 0.163 ;
      END
   END n_57645

   PIN n_57647
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.394 0.0 25.422 0.163 ;
      END
   END n_57647

   PIN n_57653
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.722 0.0 20.75 0.163 ;
      END
   END n_57653

   PIN n_58064
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 23.154 53.376 23.182 ;
      END
   END n_58064

   PIN n_58080
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.442 0.0 3.47 0.163 ;
      END
   END n_58080

   PIN n_58240
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 61.426 0.163 61.454 ;
      END
   END n_58240

   PIN n_58241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 54.77 0.163 54.798 ;
      END
   END n_58241

   PIN n_58283
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.738 0.0 34.766 0.163 ;
      END
   END n_58283

   PIN n_58284
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.954 0.0 35.982 0.163 ;
      END
   END n_58284

   PIN n_58286
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.818 76.637 32.846 76.8 ;
      END
   END n_58286

   PIN n_58527
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 43.058 53.376 43.086 ;
      END
   END n_58527

   PIN n_58659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.578 0.0 38.606 0.163 ;
      END
   END n_58659

   PIN n_58718
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.818 76.637 40.846 76.8 ;
      END
   END n_58718

   PIN n_58790
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.218 0.0 7.246 0.163 ;
      END
   END n_58790

   PIN n_58825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.458 0.163 57.486 ;
      END
   END n_58825

   PIN n_60890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 64.818 53.376 64.846 ;
      END
   END n_60890

   PIN n_61607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.082 0.163 52.11 ;
      END
   END n_61607

   PIN n_61644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.066 0.163 38.094 ;
      END
   END n_61644

   PIN n_61668
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.57 0.163 51.598 ;
      END
   END n_61668

   PIN n_6483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.018 76.637 12.046 76.8 ;
      END
   END n_6483

   PIN n_65339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 61.042 53.376 61.07 ;
      END
   END n_65339

   PIN n_67179
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 72.114 53.376 72.142 ;
      END
   END n_67179

   PIN n_7530
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.338 0.163 68.366 ;
      END
   END n_7530

   PIN n_7532
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.354 0.163 66.382 ;
      END
   END n_7532

   PIN n_7534
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.146 0.163 68.174 ;
      END
   END n_7534

   PIN n_7535
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.602 0.163 71.63 ;
      END
   END n_7535

   PIN n_7538
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.994 0.163 75.022 ;
      END
   END n_7538

   PIN n_8012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.89 0.163 75.918 ;
      END
   END n_8012

   PIN n_8483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.186 76.637 35.214 76.8 ;
      END
   END n_8483

   PIN sub_14999_49_n_82
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.546 0.163 18.574 ;
      END
   END sub_14999_49_n_82

   PIN sub_15028_54_n_56
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.762 0.163 43.79 ;
      END
   END sub_15028_54_n_56

   PIN sub_15040_54_n_63
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.202 0.163 25.23 ;
      END
   END sub_15040_54_n_63

   PIN ternarymux_ln49_0_unr5_z_7__4471875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.05 0.163 72.078 ;
      END
   END ternarymux_ln49_0_unr5_z_7__4471875

   PIN ternarymux_ln49_0_unr7_z_3__4472243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 64.69 53.376 64.718 ;
      END
   END ternarymux_ln49_0_unr7_z_3__4472243

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 53.376 76.8 ;
      LAYER V1 ;
         RECT 0.0 0.0 53.376 76.8 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 53.376 76.8 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 53.376 76.8 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 53.376 76.8 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 53.376 76.8 ;
      LAYER M1 ;
         RECT 0.0 0.0 53.376 76.8 ;
   END
END h4_mgc_edit_dist_a

MACRO h5_mgc_edit_dist_a
   CLASS BLOCK ;
   FOREIGN h5 ;
   ORIGIN 0 0 ;
   SIZE 53.376 BY 33.92 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN37857_n_42354
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.33 0.163 25.358 ;
      END
   END FE_OFN37857_n_42354

   PIN FE_OFN38247_n_35860
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 21.17 53.376 21.198 ;
      END
   END FE_OFN38247_n_35860

   PIN FE_OFN38253_n_35857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 17.97 53.376 17.998 ;
      END
   END FE_OFN38253_n_35857

   PIN FE_OFN52040_n_35867
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 25.202 53.376 25.23 ;
      END
   END FE_OFN52040_n_35867

   PIN FE_OFN52045_n_35865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 20.786 53.376 20.814 ;
      END
   END FE_OFN52045_n_35865

   PIN FE_OFN52558_n_35866
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 15.154 53.376 15.182 ;
      END
   END FE_OFN52558_n_35866

   PIN FE_OFN53041_n_35859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 21.042 53.376 21.07 ;
      END
   END FE_OFN53041_n_35859

   PIN FE_OFN53042_n_35859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 25.266 53.376 25.294 ;
      END
   END FE_OFN53042_n_35859

   PIN FE_OFN54030_n_50641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 9.202 53.376 9.23 ;
      END
   END FE_OFN54030_n_50641

   PIN FE_OFN54849_n_35866
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 21.234 53.376 21.262 ;
      END
   END FE_OFN54849_n_35866

   PIN FE_OFN69501_n_50570
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 27.058 53.376 27.086 ;
      END
   END FE_OFN69501_n_50570

   PIN FE_OFN69852_n_50569
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 27.122 53.376 27.15 ;
      END
   END FE_OFN69852_n_50569

   PIN FE_OFN72698_n_34489
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.266 33.757 1.294 33.92 ;
      END
   END FE_OFN72698_n_34489

   PIN FE_OFN87330_n_42357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.066 33.757 14.094 33.92 ;
      END
   END FE_OFN87330_n_42357

   PIN FE_OFN87336_n_42354
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.994 0.082 27.022 ;
      END
   END FE_OFN87336_n_42354

   PIN FE_OFN89085_n_34489
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.682 0.163 13.71 ;
      END
   END FE_OFN89085_n_34489

   PIN FE_OFN89086_n_34489
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.522 0.163 17.55 ;
      END
   END FE_OFN89086_n_34489

   PIN FE_OFN90160_n_57651
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.506 33.757 19.534 33.92 ;
      END
   END FE_OFN90160_n_57651

   PIN FE_OFN97083_n_50558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 21.49 53.376 21.518 ;
      END
   END FE_OFN97083_n_50558

   PIN FE_RN_1854_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 12.402 53.376 12.43 ;
      END
   END FE_RN_1854_0

   PIN FE_RN_2772_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 26.994 53.376 27.022 ;
      END
   END FE_RN_2772_0

   PIN n_35857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 20.914 53.376 20.942 ;
      END
   END n_35857

   PIN n_35859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 19.698 53.376 19.726 ;
      END
   END n_35859

   PIN n_35860
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 23.858 53.376 23.886 ;
      END
   END n_35860

   PIN n_35861
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 14.834 53.376 14.862 ;
      END
   END n_35861

   PIN n_42357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.026 0.163 31.054 ;
      END
   END n_42357

   PIN n_49961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.666 33.757 15.694 33.92 ;
      END
   END n_49961

   PIN n_49962
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.21 33.757 12.238 33.92 ;
      END
   END n_49962

   PIN n_50542
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 27.186 53.376 27.214 ;
      END
   END n_50542

   PIN n_50543
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.41 53.376 31.438 ;
      END
   END n_50543

   PIN n_50544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 27.25 53.376 27.278 ;
      END
   END n_50544

   PIN n_50552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 14.642 53.376 14.67 ;
      END
   END n_50552

   PIN n_50559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 27.314 53.376 27.342 ;
      END
   END n_50559

   PIN n_50561
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 23.986 53.376 24.014 ;
      END
   END n_50561

   PIN n_50565
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.282 53.376 31.31 ;
      END
   END n_50565

   PIN n_50566
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 27.378 53.376 27.406 ;
      END
   END n_50566

   PIN n_50571
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.346 53.376 31.374 ;
      END
   END n_50571

   PIN n_50588
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 27.442 53.376 27.47 ;
      END
   END n_50588

   PIN n_50664
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.154 53.376 31.182 ;
      END
   END n_50664

   PIN n_50670
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.65 33.757 17.678 33.92 ;
      END
   END n_50670

   PIN n_50675
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 13.682 53.376 13.71 ;
      END
   END n_50675

   PIN n_50676
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 8.69 53.376 8.718 ;
      END
   END n_50676

   PIN n_50685
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 3.058 53.376 3.086 ;
      END
   END n_50685

   PIN n_50688
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.026 33.757 47.054 33.92 ;
      END
   END n_50688

   PIN n_50692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 3.122 53.376 3.15 ;
      END
   END n_50692

   PIN n_50693
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.714 33.757 25.742 33.92 ;
      END
   END n_50693

   PIN n_50695
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.442 33.757 43.47 33.92 ;
      END
   END n_50695

   PIN n_50696
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.682 33.757 5.71 33.92 ;
      END
   END n_50696

   PIN n_50698
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.61 33.757 26.638 33.92 ;
      END
   END n_50698

   PIN n_50699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 20.146 53.376 20.174 ;
      END
   END n_50699

   PIN n_50700
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.25 33.757 51.278 33.92 ;
      END
   END n_50700

   PIN n_50701
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 3.186 53.376 3.214 ;
      END
   END n_50701

   PIN n_50702
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.682 33.757 29.71 33.92 ;
      END
   END n_50702

   PIN n_50703
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.002 33.757 30.03 33.92 ;
      END
   END n_50703

   PIN n_50704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.138 33.757 17.166 33.92 ;
      END
   END n_50704

   PIN n_50705
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 8.754 53.376 8.782 ;
      END
   END n_50705

   PIN n_50706
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 3.25 53.376 3.278 ;
      END
   END n_50706

   PIN n_50708
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.298 33.757 21.326 33.92 ;
      END
   END n_50708

   PIN n_50709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.098 33.757 34.126 33.92 ;
      END
   END n_50709

   PIN n_50711
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 14.706 53.376 14.734 ;
      END
   END n_50711

   PIN n_50712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.09 33.757 7.118 33.92 ;
      END
   END n_50712

   PIN n_52622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.698 33.757 51.726 33.92 ;
      END
   END n_52622

   PIN n_52631
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.314 33.757 3.342 33.92 ;
      END
   END n_52631

   PIN n_52632
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.218 33.757 39.246 33.92 ;
      END
   END n_52632

   PIN n_52633
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.186 33.757 35.214 33.92 ;
      END
   END n_52633

   PIN n_52634
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.346 33.757 15.374 33.92 ;
      END
   END n_52634

   PIN n_52635
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.266 33.757 41.294 33.92 ;
      END
   END n_52635

   PIN n_52639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.506 33.757 43.534 33.92 ;
      END
   END n_52639

   PIN n_52641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.45 33.757 38.478 33.92 ;
      END
   END n_52641

   PIN n_52661
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.306 33.757 24.334 33.92 ;
      END
   END n_52661

   PIN n_62553
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.258 33.757 6.286 33.92 ;
      END
   END n_62553

   PIN n_62555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.21 33.757 20.238 33.92 ;
      END
   END n_62555

   PIN n_62557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 25.458 53.376 25.486 ;
      END
   END n_62557

   PIN n_62559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.098 33.757 2.126 33.92 ;
      END
   END n_62559

   PIN n_62567
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.498 33.757 32.526 33.92 ;
      END
   END n_62567

   PIN n_62579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.202 33.757 9.23 33.92 ;
      END
   END n_62579

   PIN n_62581
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.906 33.757 9.934 33.92 ;
      END
   END n_62581

   PIN n_62582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.29 33.757 26.318 33.92 ;
      END
   END n_62582

   PIN FE_OFN49462_n_35858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 18.162 53.376 18.19 ;
      END
   END FE_OFN49462_n_35858

   PIN FE_OFN49464_n_35858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 14.962 53.376 14.99 ;
      END
   END FE_OFN49464_n_35858

   PIN FE_OFN49465_n_35858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 8.562 53.376 8.59 ;
      END
   END FE_OFN49465_n_35858

   PIN FE_OFN49995_n_42354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.714 33.757 17.742 33.92 ;
      END
   END FE_OFN49995_n_42354

   PIN FE_OFN52037_n_35867
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 14.322 53.376 14.35 ;
      END
   END FE_OFN52037_n_35867

   PIN FE_OFN52042_n_35865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 15.09 53.376 15.118 ;
      END
   END FE_OFN52042_n_35865

   PIN FE_OFN52416_n_35863
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 2.93 53.376 2.958 ;
      END
   END FE_OFN52416_n_35863

   PIN FE_OFN52418_n_35863
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 19.57 53.376 19.598 ;
      END
   END FE_OFN52418_n_35863

   PIN FE_OFN54846_n_35866
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 21.106 53.376 21.134 ;
      END
   END FE_OFN54846_n_35866

   PIN FE_OFN69978_n_46751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.202 0.163 25.23 ;
      END
   END FE_OFN69978_n_46751

   PIN FE_OFN79654_n_47488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.17 33.757 37.198 33.92 ;
      END
   END FE_OFN79654_n_47488

   PIN FE_OFN87240_n_42521
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 27.506 53.376 27.534 ;
      END
   END FE_OFN87240_n_42521

   PIN FE_OFN87249_n_35860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 21.426 53.376 21.454 ;
      END
   END FE_OFN87249_n_35860

   PIN FE_OFN87331_n_42357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.13 33.757 14.158 33.92 ;
      END
   END FE_OFN87331_n_42357

   PIN FE_OFN90096_n_47429
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.81 0.0 37.838 0.163 ;
      END
   END FE_OFN90096_n_47429

   PIN FE_OFN90159_n_57651
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.226 33.757 34.254 33.92 ;
      END
   END FE_OFN90159_n_57651

   PIN FE_OFN95252_n_47584
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.962 0.163 30.99 ;
      END
   END FE_OFN95252_n_47584

   PIN FE_RN_1856_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 12.53 53.376 12.558 ;
      END
   END FE_RN_1856_0

   PIN FE_RN_5578_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 20.082 53.376 20.11 ;
      END
   END FE_RN_5578_0

   PIN n_34489
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.218 0.163 7.246 ;
      END
   END n_34489

   PIN n_35863
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 2.802 53.376 2.83 ;
      END
   END n_35863

   PIN n_35865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 14.45 53.376 14.478 ;
      END
   END n_35865

   PIN n_42516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 25.074 53.376 25.102 ;
      END
   END n_42516

   PIN n_42517
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 19.25 53.376 19.278 ;
      END
   END n_42517

   PIN n_42518
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 30.834 53.376 30.862 ;
      END
   END n_42518

   PIN n_42520
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.09 53.376 31.118 ;
      END
   END n_42520

   PIN n_42522
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.294 30.962 53.376 30.99 ;
      END
   END n_42522

   PIN n_46750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.122 0.163 27.15 ;
      END
   END n_46750

   PIN n_46752
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.986 0.163 24.014 ;
      END
   END n_46752

   PIN n_46753
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.234 0.163 21.262 ;
      END
   END n_46753

   PIN n_47344
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.05 0.163 8.078 ;
      END
   END n_47344

   PIN n_47346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.474 0.163 15.502 ;
      END
   END n_47346

   PIN n_47348
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.41 0.163 15.438 ;
      END
   END n_47348

   PIN n_47357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 21.362 53.376 21.39 ;
      END
   END n_47357

   PIN n_47360
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 25.394 53.376 25.422 ;
      END
   END n_47360

   PIN n_47361
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.994 0.163 3.022 ;
      END
   END n_47361

   PIN n_47365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.714 0.163 9.742 ;
      END
   END n_47365

   PIN n_47366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.266 0.163 25.294 ;
      END
   END n_47366

   PIN n_47369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.386 0.163 14.414 ;
      END
   END n_47369

   PIN n_47370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 19.506 53.376 19.534 ;
      END
   END n_47370

   PIN n_47371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.154 0.163 7.182 ;
      END
   END n_47371

   PIN n_47372
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.058 0.163 3.086 ;
      END
   END n_47372

   PIN n_47373
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.986 0.163 8.014 ;
      END
   END n_47373

   PIN n_47374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.57 0.163 19.598 ;
      END
   END n_47374

   PIN n_47375
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.09 0.163 7.118 ;
      END
   END n_47375

   PIN n_47376
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.69 0.163 8.718 ;
      END
   END n_47376

   PIN n_47377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.626 0.163 8.654 ;
      END
   END n_47377

   PIN n_47378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.346 0.163 15.374 ;
      END
   END n_47378

   PIN n_47379
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.594 0.163 12.622 ;
      END
   END n_47379

   PIN n_47380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.93 0.163 2.958 ;
      END
   END n_47380

   PIN n_47383
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.506 0.163 19.534 ;
      END
   END n_47383

   PIN n_47384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.722 0.163 12.75 ;
      END
   END n_47384

   PIN n_47385
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.298 0.163 21.326 ;
      END
   END n_47385

   PIN n_47386
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.05 0.163 24.078 ;
      END
   END n_47386

   PIN n_47389
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.65 0.163 9.678 ;
      END
   END n_47389

   PIN n_47390
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.322 0.163 14.35 ;
      END
   END n_47390

   PIN n_47391
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.026 0.163 7.054 ;
      END
   END n_47391

   PIN n_47416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.962 0.163 14.99 ;
      END
   END n_47416

   PIN n_47419
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.962 0.163 14.99 ;
      END
   END n_47419

   PIN n_47427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.898 0.163 6.926 ;
      END
   END n_47427

   PIN n_47431
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.586 0.163 9.614 ;
      END
   END n_47431

   PIN n_47437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 14.578 53.376 14.606 ;
      END
   END n_47437

   PIN n_47438
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 14.514 53.376 14.542 ;
      END
   END n_47438

   PIN n_47441
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.53 0.163 12.558 ;
      END
   END n_47441

   PIN n_47442
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.658 0.163 12.686 ;
      END
   END n_47442

   PIN n_47445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.962 0.163 6.99 ;
      END
   END n_47445

   PIN n_47472
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.954 0.163 3.982 ;
      END
   END n_47472

   PIN n_47489
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.562 0.163 8.59 ;
      END
   END n_47489

   PIN n_47507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.442 0.163 19.47 ;
      END
   END n_47507

   PIN n_47510
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.226 0.163 18.254 ;
      END
   END n_47510

   PIN n_47557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.834 0.163 6.862 ;
      END
   END n_47557

   PIN n_47573
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.466 0.163 12.494 ;
      END
   END n_47573

   PIN n_47577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.866 0.163 2.894 ;
      END
   END n_47577

   PIN n_47580
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.922 0.163 7.95 ;
      END
   END n_47580

   PIN n_47581
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.802 0.163 2.83 ;
      END
   END n_47581

   PIN n_47587
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.538 33.757 47.566 33.92 ;
      END
   END n_47587

   PIN n_47589
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 21.298 53.376 21.326 ;
      END
   END n_47589

   PIN n_47591
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 31.218 53.376 31.246 ;
      END
   END n_47591

   PIN n_50557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 8.626 53.376 8.654 ;
      END
   END n_50557

   PIN n_50558
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 15.026 53.376 15.054 ;
      END
   END n_50558

   PIN n_50569
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 18.098 53.376 18.126 ;
      END
   END n_50569

   PIN n_50589
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 19.442 53.376 19.47 ;
      END
   END n_50589

   PIN n_50591
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 15.218 53.376 15.246 ;
      END
   END n_50591

   PIN n_50662
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 19.378 53.376 19.406 ;
      END
   END n_50662

   PIN n_50667
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 53.213 25.33 53.376 25.358 ;
      END
   END n_50667

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 53.376 33.92 ;
      LAYER V1 ;
         RECT 0.0 0.0 53.376 33.92 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 53.376 33.92 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 53.376 33.92 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 53.376 33.92 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 53.376 33.92 ;
      LAYER M1 ;
         RECT 0.0 0.0 53.376 33.92 ;
   END
END h5_mgc_edit_dist_a

MACRO h6_mgc_edit_dist_a
   CLASS BLOCK ;
   FOREIGN h6 ;
   ORIGIN 0 0 ;
   SIZE 51.648 BY 59.52 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN58665_n_40293
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.474 59.357 7.502 59.52 ;
      END
   END FE_OCPN58665_n_40293

   PIN FE_OCPN58699_n_40977
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.578 0.163 30.606 ;
      END
   END FE_OCPN58699_n_40977

   PIN FE_OCPN59731_n_40871
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.642 0.163 30.67 ;
      END
   END FE_OCPN59731_n_40871

   PIN FE_OCPN59829_FE_OFN27411_n_40407
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 45.234 51.648 45.262 ;
      END
   END FE_OCPN59829_FE_OFN27411_n_40407

   PIN FE_OCPN60004_n_40991
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.234 0.163 29.262 ;
      END
   END FE_OCPN60004_n_40991

   PIN FE_OCPN60013_n_40453
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.794 59.357 47.822 59.52 ;
      END
   END FE_OCPN60013_n_40453

   PIN FE_OCPN60445_n_40884
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.938 0.163 29.966 ;
      END
   END FE_OCPN60445_n_40884

   PIN FE_OCPN60817_FE_OFN50247_n_40462
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 24.626 51.648 24.654 ;
      END
   END FE_OCPN60817_FE_OFN50247_n_40462

   PIN FE_OCPN60825_n_40739
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.226 0.163 34.254 ;
      END
   END FE_OCPN60825_n_40739

   PIN FE_OCPN60829_n_40773
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 43.122 51.648 43.15 ;
      END
   END FE_OCPN60829_n_40773

   PIN FE_OCPN60889_n_40624
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 30.834 51.648 30.862 ;
      END
   END FE_OCPN60889_n_40624

   PIN FE_OCPN60892_n_40626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 29.682 51.648 29.71 ;
      END
   END FE_OCPN60892_n_40626

   PIN FE_OCPN60896_n_40916
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.218 0.163 39.246 ;
      END
   END FE_OCPN60896_n_40916

   PIN FE_OCPN61157_n_40452
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.322 0.163 30.35 ;
      END
   END FE_OCPN61157_n_40452

   PIN FE_OCPN61165_n_40736
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.722 0.163 36.75 ;
      END
   END FE_OCPN61165_n_40736

   PIN FE_OCPN61186_n_40442
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 30.77 51.648 30.798 ;
      END
   END FE_OCPN61186_n_40442

   PIN FE_OCPN61190_n_40385
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.33 0.163 33.358 ;
      END
   END FE_OCPN61190_n_40385

   PIN FE_OCPN61194_n_40543
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.386 0.163 30.414 ;
      END
   END FE_OCPN61194_n_40543

   PIN FE_OCPN61198_FE_OFN4340_n_40574
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.682 59.357 21.71 59.52 ;
      END
   END FE_OCPN61198_FE_OFN4340_n_40574

   PIN FE_OCPN61200_FE_OFN26050_n_40461
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 48.114 51.648 48.142 ;
      END
   END FE_OCPN61200_FE_OFN26050_n_40461

   PIN FE_OCPN61205_n_40748
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.706 0.163 30.734 ;
      END
   END FE_OCPN61205_n_40748

   PIN FE_OCPN61340_n_40638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.274 59.357 36.302 59.52 ;
      END
   END FE_OCPN61340_n_40638

   PIN FE_OCPN61708_n_40671
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.002 0.163 54.03 ;
      END
   END FE_OCPN61708_n_40671

   PIN FE_OCPN62299_FE_OFN53822_n_40455
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.594 0.163 36.622 ;
      END
   END FE_OCPN62299_FE_OFN53822_n_40455

   PIN FE_OCPN62464_n_40460
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.402 0.163 20.43 ;
      END
   END FE_OCPN62464_n_40460

   PIN FE_OCPN62757_n_40522
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.986 0.163 48.014 ;
      END
   END FE_OCPN62757_n_40522

   PIN FE_OCPN62762_n_40389
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 52.082 51.648 52.11 ;
      END
   END FE_OCPN62762_n_40389

   PIN FE_OCPN62778_n_40539
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.682 0.163 53.71 ;
      END
   END FE_OCPN62778_n_40539

   PIN FE_OCPN63314_n_40689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.378 0.163 11.406 ;
      END
   END FE_OCPN63314_n_40689

   PIN FE_OCPN63402_n_40695
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.626 59.357 24.654 59.52 ;
      END
   END FE_OCPN63402_n_40695

   PIN FE_OCPN63686_n_40655
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.81 59.357 21.838 59.52 ;
      END
   END FE_OCPN63686_n_40655

   PIN FE_OCPN63879_n_40667
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.05 59.357 32.078 59.52 ;
      END
   END FE_OCPN63879_n_40667

   PIN FE_OCPN76175_n_40685
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.162 59.357 10.19 59.52 ;
      END
   END FE_OCPN76175_n_40685

   PIN FE_OCPN76176_n_40685
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.034 59.357 42.062 59.52 ;
      END
   END FE_OCPN76176_n_40685

   PIN FE_OCPN76225_n_40728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.794 0.163 15.822 ;
      END
   END FE_OCPN76225_n_40728

   PIN FE_OCPN76871_n_40344
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.786 0.163 44.814 ;
      END
   END FE_OCPN76871_n_40344

   PIN FE_OCPN76899_n_40732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.706 0.163 6.734 ;
      END
   END FE_OCPN76899_n_40732

   PIN FE_OCPN77057_n_40646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.658 0.163 20.686 ;
      END
   END FE_OCPN77057_n_40646

   PIN FE_OCPN77058_n_40646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.754 0.163 24.782 ;
      END
   END FE_OCPN77058_n_40646

   PIN FE_OCPN78169_n_40634
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.33 59.357 33.358 59.52 ;
      END
   END FE_OCPN78169_n_40634

   PIN FE_OCPN78237_FE_OFN3733_n_40730
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.178 0.163 16.206 ;
      END
   END FE_OCPN78237_FE_OFN3733_n_40730

   PIN FE_OCPN95535_n_40744
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 42.29 51.648 42.318 ;
      END
   END FE_OCPN95535_n_40744

   PIN FE_OCPN95538_FE_OFN90000_n_40684
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.994 0.163 19.022 ;
      END
   END FE_OCPN95538_FE_OFN90000_n_40684

   PIN FE_OCPN95613_FE_OFN89862_n_40309
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 39.346 51.648 39.374 ;
      END
   END FE_OCPN95613_FE_OFN89862_n_40309

   PIN FE_OCPN95619_n_40607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 47.602 51.648 47.63 ;
      END
   END FE_OCPN95619_n_40607

   PIN FE_OCPN95761_n_40465
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.09 59.357 39.118 59.52 ;
      END
   END FE_OCPN95761_n_40465

   PIN FE_OCPN95853_FE_OFN90041_n_40381
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 51.485 57.202 51.648 57.23 ;
      END
   END FE_OCPN95853_FE_OFN90041_n_40381

   PIN FE_OCP_DRV_N76452_FE_OFN67430_n_40505
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.634 0.163 27.662 ;
      END
   END FE_OCP_DRV_N76452_FE_OFN67430_n_40505

   PIN FE_OCP_DRV_N76464_FE_OFN66917_n_40672
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 45.298 51.648 45.326 ;
      END
   END FE_OCP_DRV_N76464_FE_OFN66917_n_40672

   PIN FE_OCP_DRV_N78200_FE_OFN37047_n_35919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.186 0.163 11.214 ;
      END
   END FE_OCP_DRV_N78200_FE_OFN37047_n_35919

   PIN FE_OFN3336_n_57614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.97 59.357 1.998 59.52 ;
      END
   END FE_OFN3336_n_57614

   PIN FE_OFN35849_n_52031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.122 59.357 19.15 59.52 ;
      END
   END FE_OFN35849_n_52031

   PIN FE_OFN35858_n_52027
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.322 59.357 22.35 59.52 ;
      END
   END FE_OFN35858_n_52027

   PIN FE_OFN35873_n_52030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.106 59.357 13.134 59.52 ;
      END
   END FE_OFN35873_n_52030

   PIN FE_OFN35875_n_52030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.85 59.357 4.878 59.52 ;
      END
   END FE_OFN35875_n_52030

   PIN FE_OFN35909_n_52083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.49 0.163 13.518 ;
      END
   END FE_OFN35909_n_52083

   PIN FE_OFN35925_n_52086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 20.082 0.163 20.11 ;
      END
   END FE_OFN35925_n_52086

   PIN FE_OFN35933_n_52028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.018 59.357 36.046 59.52 ;
      END
   END FE_OFN35933_n_52028

   PIN FE_OFN35937_n_52028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.426 59.438 5.454 59.52 ;
      END
   END FE_OFN35937_n_52028

   PIN FE_OFN36907_n_35904
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.602 0.163 47.63 ;
      END
   END FE_OFN36907_n_35904

   PIN FE_OFN36908_n_35904
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.122 59.438 19.15 59.52 ;
      END
   END FE_OFN36908_n_35904

   PIN FE_OFN36982_n_45345
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.362 59.357 13.39 59.52 ;
      END
   END FE_OFN36982_n_45345

   PIN FE_OFN37047_n_35919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.298 0.163 13.326 ;
      END
   END FE_OFN37047_n_35919

   PIN FE_OFN4914_n_56419
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.298 0.163 45.326 ;
      END
   END FE_OFN4914_n_56419

   PIN FE_OFN50279_n_52028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.562 0.163 24.59 ;
      END
   END FE_OFN50279_n_52028

   PIN FE_OFN50280_n_52028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.354 0.163 42.382 ;
      END
   END FE_OFN50280_n_52028

   PIN FE_OFN50334_n_52030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.186 59.357 19.214 59.52 ;
      END
   END FE_OFN50334_n_52030

   PIN FE_OFN50335_n_52030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.506 0.163 27.534 ;
      END
   END FE_OFN50335_n_52030

   PIN FE_OFN53021_n_40337
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.898 0.163 38.926 ;
      END
   END FE_OFN53021_n_40337

   PIN FE_OFN53588_n_40797
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 19.314 51.648 19.342 ;
      END
   END FE_OFN53588_n_40797

   PIN FE_OFN53589_n_40797
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.258 0.163 22.286 ;
      END
   END FE_OFN53589_n_40797

   PIN FE_OFN53785_n_52084
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.05 0.163 16.078 ;
      END
   END FE_OFN53785_n_52084

   PIN FE_OFN53787_n_52080
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.626 59.357 8.654 59.52 ;
      END
   END FE_OFN53787_n_52080

   PIN FE_OFN53788_n_52080
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.362 0.163 45.39 ;
      END
   END FE_OFN53788_n_52080

   PIN FE_OFN53789_n_52080
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.914 59.357 12.942 59.52 ;
      END
   END FE_OFN53789_n_52080

   PIN FE_OFN53790_n_52080
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.898 0.163 30.926 ;
      END
   END FE_OFN53790_n_52080

   PIN FE_OFN53791_n_52027
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.938 0.163 13.966 ;
      END
   END FE_OFN53791_n_52027

   PIN FE_OFN53792_n_52027
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.754 59.357 24.782 59.52 ;
      END
   END FE_OFN53792_n_52027

   PIN FE_OFN53795_n_52027
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.426 59.357 13.454 59.52 ;
      END
   END FE_OFN53795_n_52027

   PIN FE_OFN53796_n_52087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.442 0.163 27.47 ;
      END
   END FE_OFN53796_n_52087

   PIN FE_OFN53797_n_52087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.298 59.438 13.326 59.52 ;
      END
   END FE_OFN53797_n_52087

   PIN FE_OFN53798_n_52087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.17 59.357 13.198 59.52 ;
      END
   END FE_OFN53798_n_52087

   PIN FE_OFN53806_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.682 59.357 5.71 59.52 ;
      END
   END FE_OFN53806_n_52029

   PIN FE_OFN53807_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.842 0.163 33.87 ;
      END
   END FE_OFN53807_n_52029

   PIN FE_OFN53808_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.882 59.438 24.91 59.52 ;
      END
   END FE_OFN53808_n_52029

   PIN FE_OFN53810_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.386 59.357 38.414 59.52 ;
      END
   END FE_OFN53810_n_52029

   PIN FE_OFN53813_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.29 0.163 34.318 ;
      END
   END FE_OFN53813_n_52029

   PIN FE_OFN53847_n_52031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.482 59.357 10.51 59.52 ;
      END
   END FE_OFN53847_n_52031

   PIN FE_OFN53848_n_52031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.082 0.163 20.11 ;
      END
   END FE_OFN53848_n_52031

   PIN FE_OFN53852_n_52081
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.874 0.163 53.902 ;
      END
   END FE_OFN53852_n_52081

   PIN FE_OFN53929_n_52024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.554 0.163 45.582 ;
      END
   END FE_OFN53929_n_52024

   PIN FE_OFN53930_n_52024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.722 59.357 4.75 59.52 ;
      END
   END FE_OFN53930_n_52024

   PIN FE_OFN53951_n_40618
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 24.562 51.648 24.59 ;
      END
   END FE_OFN53951_n_40618

   PIN FE_OFN53970_n_40476
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.858 0.163 15.886 ;
      END
   END FE_OFN53970_n_40476

   PIN FE_OFN53975_n_52082
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.002 0.163 30.03 ;
      END
   END FE_OFN53975_n_52082

   PIN FE_OFN53976_n_52082
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.282 0.163 39.31 ;
      END
   END FE_OFN53976_n_52082

   PIN FE_OFN54053_n_53997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.418 0.163 2.446 ;
      END
   END FE_OFN54053_n_53997

   PIN FE_OFN55531_n_45338
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.354 59.357 10.382 59.52 ;
      END
   END FE_OFN55531_n_45338

   PIN FE_OFN55721_n_52025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.394 59.357 41.422 59.52 ;
      END
   END FE_OFN55721_n_52025

   PIN FE_OFN55722_n_52025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.882 0.163 24.91 ;
      END
   END FE_OFN55722_n_52025

   PIN FE_OFN55723_n_52025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.738 0.163 50.766 ;
      END
   END FE_OFN55723_n_52025

   PIN FE_OFN55724_n_52025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.922 59.357 15.95 59.52 ;
      END
   END FE_OFN55724_n_52025

   PIN FE_OFN55763_n_52086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.41 59.357 7.438 59.52 ;
      END
   END FE_OFN55763_n_52086

   PIN FE_OFN55765_n_52086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.994 59.438 19.022 59.52 ;
      END
   END FE_OFN55765_n_52086

   PIN FE_OFN55829_n_52085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.098 59.357 2.126 59.52 ;
      END
   END FE_OFN55829_n_52085

   PIN FE_OFN55830_n_52085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.49 59.357 13.518 59.52 ;
      END
   END FE_OFN55830_n_52085

   PIN FE_OFN55832_n_52085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.498 0.163 16.526 ;
      END
   END FE_OFN55832_n_52085

   PIN FE_OFN64709_n_40441
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.858 59.357 47.886 59.52 ;
      END
   END FE_OFN64709_n_40441

   PIN FE_OFN64798_n_40578
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.362 59.357 21.39 59.52 ;
      END
   END FE_OFN64798_n_40578

   PIN FE_OFN64923_n_40587
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.69 59.357 24.718 59.52 ;
      END
   END FE_OFN64923_n_40587

   PIN FE_OFN67632_n_40380
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.322 0.163 22.35 ;
      END
   END FE_OFN67632_n_40380

   PIN FE_OFN67675_n_41246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.362 0.163 13.39 ;
      END
   END FE_OFN67675_n_41246

   PIN FE_OFN68512_n_40584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.866 59.357 18.894 59.52 ;
      END
   END FE_OFN68512_n_40584

   PIN FE_OFN68513_n_40584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.466 0.163 20.494 ;
      END
   END FE_OFN68513_n_40584

   PIN FE_OFN68659_n_41001
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.818 0.163 56.846 ;
      END
   END FE_OFN68659_n_41001

   PIN FE_OFN68752_n_40468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.93 59.357 18.958 59.52 ;
      END
   END FE_OFN68752_n_40468

   PIN FE_OFN69011_n_40742
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 43.186 51.648 43.214 ;
      END
   END FE_OFN69011_n_40742

   PIN FE_OFN69206_n_40725
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.81 0.163 21.838 ;
      END
   END FE_OFN69206_n_40725

   PIN FE_OFN69664_n_40499
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.69 0.163 24.718 ;
      END
   END FE_OFN69664_n_40499

   PIN FE_OFN69889_n_40422
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.962 0.163 30.99 ;
      END
   END FE_OFN69889_n_40422

   PIN FE_OFN70042_n_40615
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.69 59.357 24.718 59.52 ;
      END
   END FE_OFN70042_n_40615

   PIN FE_OFN79586_n_40690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.05 59.357 16.078 59.52 ;
      END
   END FE_OFN79586_n_40690

   PIN FE_OFN79626_n_40616
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 51.485 50.994 51.648 51.022 ;
      END
   END FE_OFN79626_n_40616

   PIN FE_OFN80551_n_41085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 48.05 51.648 48.078 ;
      END
   END FE_OFN80551_n_41085

   PIN FE_OFN81546_n_40579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 36.594 51.648 36.622 ;
      END
   END FE_OFN81546_n_40579

   PIN FE_OFN82254_n_40562
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.85 0.163 20.878 ;
      END
   END FE_OFN82254_n_40562

   PIN FE_OFN82720_n_40745
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.93 0.163 50.958 ;
      END
   END FE_OFN82720_n_40745

   PIN FE_OFN84632_n_45520
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 53.554 51.648 53.582 ;
      END
   END FE_OFN84632_n_45520

   PIN FE_OFN89562_n_40600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.994 0.163 51.022 ;
      END
   END FE_OFN89562_n_40600

   PIN FE_OFN89690_n_40666
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 38.706 51.648 38.734 ;
      END
   END FE_OFN89690_n_40666

   PIN FE_OFN89775_n_40818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.418 0.163 42.446 ;
      END
   END FE_OFN89775_n_40818

   PIN FE_OFN89783_n_41094
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.522 0.163 25.55 ;
      END
   END FE_OFN89783_n_41094

   PIN FE_OFN89834_n_40765
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.026 59.357 7.054 59.52 ;
      END
   END FE_OFN89834_n_40765

   PIN FE_OFN89889_n_40579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 25.01 51.648 25.038 ;
      END
   END FE_OFN89889_n_40579

   PIN FE_OFN89896_n_40690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.45 59.357 30.478 59.52 ;
      END
   END FE_OFN89896_n_40690

   PIN FE_OFN89931_n_41129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.41 59.357 39.438 59.52 ;
      END
   END FE_OFN89931_n_41129

   PIN FE_OFN89946_n_40368
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.386 0.163 22.414 ;
      END
   END FE_OFN89946_n_40368

   PIN FE_OFN89969_n_40791
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.37 59.357 48.398 59.52 ;
      END
   END FE_OFN89969_n_40791

   PIN FE_OFN89991_n_40449
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.554 0.163 13.582 ;
      END
   END FE_OFN89991_n_40449

   PIN FE_OFN89995_n_40526
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.098 59.357 42.126 59.52 ;
      END
   END FE_OFN89995_n_40526

   PIN FE_OFN89996_n_40526
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 38.77 51.648 38.798 ;
      END
   END FE_OFN89996_n_40526

   PIN FE_OFN90072_FE_OCPN57974_n_40531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 42.354 51.648 42.382 ;
      END
   END FE_OFN90072_FE_OCPN57974_n_40531

   PIN FE_OFN90077_n_40436
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.562 59.357 24.59 59.52 ;
      END
   END FE_OFN90077_n_40436

   PIN FE_OFN90083_n_40637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.426 0.163 45.454 ;
      END
   END FE_OFN90083_n_40637

   PIN FE_OFN92416_n_40768
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.482 0.163 42.51 ;
      END
   END FE_OFN92416_n_40768

   PIN FE_OFN92692_n_40849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.618 0.163 13.646 ;
      END
   END FE_OFN92692_n_40849

   PIN FE_OFN92693_n_40849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.682 0.163 13.71 ;
      END
   END FE_OFN92693_n_40849

   PIN FE_OFN92898_n_40770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.194 0.163 38.222 ;
      END
   END FE_OFN92898_n_40770

   PIN FE_OFN93228_n_40835
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.818 0.163 24.846 ;
      END
   END FE_OFN93228_n_40835

   PIN FE_OFN95235_n_40680
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.946 0.163 24.974 ;
      END
   END FE_OFN95235_n_40680

   PIN FE_OFN95251_n_40692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.218 59.357 31.246 59.52 ;
      END
   END FE_OFN95251_n_40692

   PIN FE_OFN95268_n_40689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.442 0.163 11.47 ;
      END
   END FE_OFN95268_n_40689

   PIN FE_OFN96061_FE_OCPN59260_n_40732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.866 0.163 18.894 ;
      END
   END FE_OFN96061_FE_OCPN59260_n_40732

   PIN FE_OFN96635_n_41231
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.658 0.163 36.686 ;
      END
   END FE_OFN96635_n_41231

   PIN FE_OFN96853_FE_OCPN61163_n_40472
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.77 0.163 30.798 ;
      END
   END FE_OFN96853_FE_OCPN61163_n_40472

   PIN FE_OFN96935_n_40586
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.306 0.163 48.334 ;
      END
   END FE_OFN96935_n_40586

   PIN FE_OFN96959_n_40592
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.57 59.357 27.598 59.52 ;
      END
   END FE_OFN96959_n_40592

   PIN FE_OFN97148_n_41111
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.906 0.163 33.934 ;
      END
   END FE_OFN97148_n_41111

   PIN FE_OFN97292_n_40798
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.634 59.357 27.662 59.52 ;
      END
   END FE_OFN97292_n_40798

   PIN FE_OFN97614_FE_OCPN61281_n_40613
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.634 59.357 27.662 59.52 ;
      END
   END FE_OFN97614_FE_OCPN61281_n_40613

   PIN FE_RN_3275_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.754 59.357 24.782 59.52 ;
      END
   END FE_RN_3275_0

   PIN FE_RN_3761_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.01 0.163 25.038 ;
      END
   END FE_RN_3761_0

   PIN FE_RN_541_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.97 59.357 9.998 59.52 ;
      END
   END FE_RN_541_0

   PIN n_44333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 50.994 51.648 51.022 ;
      END
   END n_44333

   PIN n_44349
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 51.058 51.648 51.086 ;
      END
   END n_44349

   PIN n_44353
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.322 59.357 6.35 59.52 ;
      END
   END n_44353

   PIN n_44354
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.914 59.357 44.942 59.52 ;
      END
   END n_44354

   PIN n_44355
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 6.642 51.648 6.67 ;
      END
   END n_44355

   PIN n_44356
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 2.162 51.648 2.19 ;
      END
   END n_44356

   PIN n_44359
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 47.666 51.648 47.694 ;
      END
   END n_44359

   PIN n_44383
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 34.226 51.648 34.254 ;
      END
   END n_44383

   PIN n_44384
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.362 59.357 37.39 59.52 ;
      END
   END n_44384

   PIN n_45336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.234 59.357 13.262 59.52 ;
      END
   END n_45336

   PIN n_45339
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.474 59.357 7.502 59.52 ;
      END
   END n_45339

   PIN n_45342
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.098 59.357 34.126 59.52 ;
      END
   END n_45342

   PIN n_45343
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.922 59.357 7.95 59.52 ;
      END
   END n_45343

   PIN n_45344
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.682 0.163 45.71 ;
      END
   END n_45344

   PIN n_45346
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.298 59.357 13.326 59.52 ;
      END
   END n_45346

   PIN n_52024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.994 59.357 19.022 59.52 ;
      END
   END n_52024

   PIN n_52082
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.946 59.357 24.974 59.52 ;
      END
   END n_52082

   PIN n_53966
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.578 0.163 22.606 ;
      END
   END n_53966

   PIN n_53968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.146 0.163 28.174 ;
      END
   END n_53968

   PIN n_53995
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.586 0.163 25.614 ;
      END
   END n_53995

   PIN n_53996
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.074 0.163 25.102 ;
      END
   END n_53996

   PIN n_54003
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.114 59.357 16.142 59.52 ;
      END
   END n_54003

   PIN n_54014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.17 59.357 13.198 59.52 ;
      END
   END n_54014

   PIN n_54043
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.434 0.163 16.462 ;
      END
   END n_54043

   PIN n_54057
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.53 0.163 20.558 ;
      END
   END n_54057

   PIN n_54098
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.314 0.163 43.342 ;
      END
   END n_54098

   PIN n_54186
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.218 59.357 7.246 59.52 ;
      END
   END n_54186

   PIN n_54198
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.786 59.357 4.814 59.52 ;
      END
   END n_54198

   PIN n_54215
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.978 59.357 5.006 59.52 ;
      END
   END n_54215

   PIN n_54238
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.282 59.357 7.31 59.52 ;
      END
   END n_54238

   PIN n_54239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.346 59.357 7.374 59.52 ;
      END
   END n_54239

   PIN n_56417
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.802 59.357 18.83 59.52 ;
      END
   END n_56417

   PIN n_56423
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.034 59.357 2.062 59.52 ;
      END
   END n_56423

   PIN n_56424
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.714 59.357 1.742 59.52 ;
      END
   END n_56424

   PIN n_56425
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 36.594 0.163 36.622 ;
      END
   END n_56425

   PIN n_56426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.346 0.163 39.374 ;
      END
   END n_56426

   PIN n_56429
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.122 0.163 11.15 ;
      END
   END n_56429

   PIN n_57591
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.882 59.357 24.91 59.52 ;
      END
   END n_57591

   PIN n_58389
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.962 0.163 38.99 ;
      END
   END n_58389

   PIN n_58593
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.778 59.357 1.806 59.52 ;
      END
   END n_58593

   PIN n_58665
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.202 0.163 57.23 ;
      END
   END n_58665

   PIN FE_OCPN57928_n_40786
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.338 0.163 20.366 ;
      END
   END FE_OCPN57928_n_40786

   PIN FE_OCPN57974_n_40531
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.026 0.163 7.054 ;
      END
   END FE_OCPN57974_n_40531

   PIN FE_OCPN58664_n_40293
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.922 0.163 15.95 ;
      END
   END FE_OCPN58664_n_40293

   PIN FE_OCPN58691_n_40304
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 19.314 0.163 19.342 ;
      END
   END FE_OCPN58691_n_40304

   PIN FE_OCPN58698_n_40977
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.37 0.163 16.398 ;
      END
   END FE_OCPN58698_n_40977

   PIN FE_OCPN59256_n_40667
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.266 0.163 57.294 ;
      END
   END FE_OCPN59256_n_40667

   PIN FE_OCPN59258_n_40370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.954 0.163 27.982 ;
      END
   END FE_OCPN59258_n_40370

   PIN FE_OCPN59262_n_40728
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.234 0.163 13.262 ;
      END
   END FE_OCPN59262_n_40728

   PIN FE_OCPN59729_n_40871
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.17 0.163 29.198 ;
      END
   END FE_OCPN59729_n_40871

   PIN FE_OCPN59744_n_40606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.354 0.163 2.382 ;
      END
   END FE_OCPN59744_n_40606

   PIN FE_OCPN59823_n_40673
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.69 59.357 16.718 59.52 ;
      END
   END FE_OCPN59823_n_40673

   PIN FE_OCPN59828_FE_OFN27411_n_40407
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.914 0.163 36.942 ;
      END
   END FE_OCPN59828_FE_OFN27411_n_40407

   PIN FE_OCPN59987_n_40388
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 23.026 0.163 23.054 ;
      END
   END FE_OCPN59987_n_40388

   PIN FE_OCPN60002_n_40991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.106 0.163 29.134 ;
      END
   END FE_OCPN60002_n_40991

   PIN FE_OCPN60011_n_40453
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.226 59.357 26.254 59.52 ;
      END
   END FE_OCPN60011_n_40453

   PIN FE_OCPN60444_n_40884
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.874 0.163 29.902 ;
      END
   END FE_OCPN60444_n_40884

   PIN FE_OCPN60815_FE_OFN50247_n_40462
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.746 0.163 29.774 ;
      END
   END FE_OCPN60815_FE_OFN50247_n_40462

   PIN FE_OCPN60824_n_40739
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.53 0.163 36.558 ;
      END
   END FE_OCPN60824_n_40739

   PIN FE_OCPN60827_n_40753
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 38.642 51.648 38.67 ;
      END
   END FE_OCPN60827_n_40753

   PIN FE_OCPN60828_n_40773
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.25 0.163 43.278 ;
      END
   END FE_OCPN60828_n_40773

   PIN FE_OCPN60887_n_40624
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.29 0.163 34.318 ;
      END
   END FE_OCPN60887_n_40624

   PIN FE_OCPN60890_n_40626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 29.682 0.163 29.71 ;
      END
   END FE_OCPN60890_n_40626

   PIN FE_OCPN60895_n_40916
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.162 0.163 34.19 ;
      END
   END FE_OCPN60895_n_40916

   PIN FE_OCPN60898_FE_OFN3733_n_40730
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.29 0.163 2.318 ;
      END
   END FE_OCPN60898_FE_OFN3733_n_40730

   PIN FE_OCPN61161_n_40733
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.114 0.163 16.142 ;
      END
   END FE_OCPN61161_n_40733

   PIN FE_OCPN61163_n_40472
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.042 0.163 29.07 ;
      END
   END FE_OCPN61163_n_40472

   PIN FE_OCPN61164_n_40736
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.65 0.163 33.678 ;
      END
   END FE_OCPN61164_n_40736

   PIN FE_OCPN61170_n_40664
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.658 59.357 4.686 59.52 ;
      END
   END FE_OCPN61170_n_40664

   PIN FE_OCPN61178_n_40494
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.266 0.163 25.294 ;
      END
   END FE_OCPN61178_n_40494

   PIN FE_OCPN61180_FE_OFN26782_n_40493
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 34.162 51.648 34.19 ;
      END
   END FE_OCPN61180_FE_OFN26782_n_40493

   PIN FE_OCPN61184_n_40665
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.618 0.163 53.646 ;
      END
   END FE_OCPN61184_n_40665

   PIN FE_OCPN61188_n_40458
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.778 0.163 33.806 ;
      END
   END FE_OCPN61188_n_40458

   PIN FE_OCPN61189_n_40385
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.73 0.163 15.758 ;
      END
   END FE_OCPN61189_n_40385

   PIN FE_OCPN61193_n_40543
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.93 0.163 18.958 ;
      END
   END FE_OCPN61193_n_40543

   PIN FE_OCPN61197_FE_OFN4340_n_40574
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.282 0.163 7.31 ;
      END
   END FE_OCPN61197_FE_OFN4340_n_40574

   PIN FE_OCPN61199_FE_OFN26050_n_40461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 43.186 0.163 43.214 ;
      END
   END FE_OCPN61199_FE_OFN26050_n_40461

   PIN FE_OCPN61202_n_40700
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.234 0.163 45.262 ;
      END
   END FE_OCPN61202_n_40700

   PIN FE_OCPN61281_n_40613
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.066 0.163 54.094 ;
      END
   END FE_OCPN61281_n_40613

   PIN FE_OCPN61334_n_40487
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.626 0.163 24.654 ;
      END
   END FE_OCPN61334_n_40487

   PIN FE_OCPN61703_n_40614
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.89 0.163 27.918 ;
      END
   END FE_OCPN61703_n_40614

   PIN FE_OCPN61705_n_40652
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.826 0.163 27.854 ;
      END
   END FE_OCPN61705_n_40652

   PIN FE_OCPN61706_n_40671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.938 0.163 53.966 ;
      END
   END FE_OCPN61706_n_40671

   PIN FE_OCPN61855_FE_OFN53951_n_40618
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 25.074 51.648 25.102 ;
      END
   END FE_OCPN61855_FE_OFN53951_n_40618

   PIN FE_OCPN61880_FE_OFN21562_n_40405
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.186 0.163 51.214 ;
      END
   END FE_OCPN61880_FE_OFN21562_n_40405

   PIN FE_OCPN61918_FE_OFN53968_n_40476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.666 0.163 15.694 ;
      END
   END FE_OCPN61918_FE_OFN53968_n_40476

   PIN FE_OCPN62235_n_40789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.81 0.163 29.838 ;
      END
   END FE_OCPN62235_n_40789

   PIN FE_OCPN62246_n_40447
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.226 0.163 2.254 ;
      END
   END FE_OCPN62246_n_40447

   PIN FE_OCPN62248_n_40471
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.29 59.357 10.318 59.52 ;
      END
   END FE_OCPN62248_n_40471

   PIN FE_OCPN62288_FE_OFN53950_n_40618
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.682 0.163 29.71 ;
      END
   END FE_OCPN62288_FE_OFN53950_n_40618

   PIN FE_OCPN62466_n_40460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.914 0.163 4.942 ;
      END
   END FE_OCPN62466_n_40460

   PIN FE_OCPN62755_n_40522
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.466 0.163 36.494 ;
      END
   END FE_OCPN62755_n_40522

   PIN FE_OCPN62760_n_40389
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.146 0.163 52.174 ;
      END
   END FE_OCPN62760_n_40389

   PIN FE_OCPN62777_n_40539
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.122 0.163 51.15 ;
      END
   END FE_OCPN62777_n_40539

   PIN FE_OCPN63398_n_41185
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.866 0.163 50.894 ;
      END
   END FE_OCPN63398_n_41185

   PIN FE_OCPN63401_n_40695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.834 0.163 38.862 ;
      END
   END FE_OCPN63401_n_40695

   PIN FE_OCPN63684_n_40655
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.962 0.163 46.99 ;
      END
   END FE_OCPN63684_n_40655

   PIN FE_OCPN63702_n_40513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.962 0.163 6.99 ;
      END
   END FE_OCPN63702_n_40513

   PIN FE_OCPN63974_n_40634
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.058 59.357 11.086 59.52 ;
      END
   END FE_OCPN63974_n_40634

   PIN FE_OCPN76163_n_40638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.146 59.357 36.174 59.52 ;
      END
   END FE_OCPN76163_n_40638

   PIN FE_OCPN76302_FE_OFN67600_n_40588
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.194 0.163 22.222 ;
      END
   END FE_OCPN76302_FE_OFN67600_n_40588

   PIN FE_OCPN76722_n_40452
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.978 0.163 5.006 ;
      END
   END FE_OCPN76722_n_40452

   PIN FE_OCPN76870_n_40344
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.274 0.163 20.302 ;
      END
   END FE_OCPN76870_n_40344

   PIN FE_OCPN77056_n_40657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.554 0.163 53.582 ;
      END
   END FE_OCPN77056_n_40657

   PIN FE_OCPN95432_FE_OFN89660_n_40792
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.402 0.163 36.43 ;
      END
   END FE_OCPN95432_FE_OFN89660_n_40792

   PIN FE_OCPN95534_n_40744
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 38.706 0.163 38.734 ;
      END
   END FE_OCPN95534_n_40744

   PIN FE_OCPN95536_FE_OFN90000_n_40684
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.634 0.163 11.662 ;
      END
   END FE_OCPN95536_FE_OFN90000_n_40684

   PIN FE_OCPN95612_FE_OFN89862_n_40309
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.618 0.163 45.646 ;
      END
   END FE_OCPN95612_FE_OFN89862_n_40309

   PIN FE_OCPN95618_n_40607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.17 0.163 45.198 ;
      END
   END FE_OCPN95618_n_40607

   PIN FE_OCPN95760_n_40465
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.034 0.163 58.062 ;
      END
   END FE_OCPN95760_n_40465

   PIN FE_OCPN99043_n_40638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.058 0.163 51.086 ;
      END
   END FE_OCPN99043_n_40638

   PIN FE_OCP_DRV_N78196_n_40785
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.298 59.357 37.326 59.52 ;
      END
   END FE_OCP_DRV_N78196_n_40785

   PIN FE_OCP_DRV_N78718_FE_OFN69107_n_40425
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.434 0.163 16.462 ;
      END
   END FE_OCP_DRV_N78718_FE_OFN69107_n_40425

   PIN FE_OCP_DRV_N99398_FE_OFN98007_n_35906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.514 59.357 30.542 59.52 ;
      END
   END FE_OCP_DRV_N99398_FE_OFN98007_n_35906

   PIN FE_OFN11400_n_40826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.37 0.163 16.398 ;
      END
   END FE_OFN11400_n_40826

   PIN FE_OFN36963_n_35917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.698 59.357 27.726 59.52 ;
      END
   END FE_OFN36963_n_35917

   PIN FE_OFN36981_n_45345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.458 59.357 25.486 59.52 ;
      END
   END FE_OFN36981_n_45345

   PIN FE_OFN37043_n_35919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.018 0.163 28.046 ;
      END
   END FE_OFN37043_n_35919

   PIN FE_OFN37045_n_35919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.458 0.163 25.486 ;
      END
   END FE_OFN37045_n_35919

   PIN FE_OFN37046_n_35919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.29 0.163 42.318 ;
      END
   END FE_OFN37046_n_35919

   PIN FE_OFN37067_n_35921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.17 0.163 13.198 ;
      END
   END FE_OFN37067_n_35921

   PIN FE_OFN46443_n_35921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.394 0.163 25.422 ;
      END
   END FE_OFN46443_n_35921

   PIN FE_OFN46639_n_35902
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.986 59.357 32.014 59.52 ;
      END
   END FE_OFN46639_n_35902

   PIN FE_OFN46654_n_35904
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.418 59.357 10.446 59.52 ;
      END
   END FE_OFN46654_n_35904

   PIN FE_OFN49989_n_40350
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 45.554 0.163 45.582 ;
      END
   END FE_OFN49989_n_40350

   PIN FE_OFN49990_n_40689
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.122 0.163 11.15 ;
      END
   END FE_OFN49990_n_40689

   PIN FE_OFN50159_n_51368
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.922 59.357 47.95 59.52 ;
      END
   END FE_OFN50159_n_51368

   PIN FE_OFN50261_n_51366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.074 59.357 49.102 59.52 ;
      END
   END FE_OFN50261_n_51366

   PIN FE_OFN50310_n_40737
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.338 0.163 36.366 ;
      END
   END FE_OFN50310_n_40737

   PIN FE_OFN52335_n_45520
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.202 59.357 49.23 59.52 ;
      END
   END FE_OFN52335_n_45520

   PIN FE_OFN5281_n_40391
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 42.354 0.163 42.382 ;
      END
   END FE_OFN5281_n_40391

   PIN FE_OFN53002_n_40279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.106 0.163 45.134 ;
      END
   END FE_OFN53002_n_40279

   PIN FE_OFN53022_n_40337
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.714 0.163 33.742 ;
      END
   END FE_OFN53022_n_40337

   PIN FE_OFN53283_n_40791
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.922 0.163 47.95 ;
      END
   END FE_OFN53283_n_40791

   PIN FE_OFN53291_n_41258
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.314 0.163 11.342 ;
      END
   END FE_OFN53291_n_41258

   PIN FE_OFN53587_n_40797
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.874 0.163 13.902 ;
      END
   END FE_OFN53587_n_40797

   PIN FE_OFN53642_n_40692
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.042 59.357 13.07 59.52 ;
      END
   END FE_OFN53642_n_40692

   PIN FE_OFN53722_n_40501
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.594 0.163 20.622 ;
      END
   END FE_OFN53722_n_40501

   PIN FE_OFN53780_n_52084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.082 59.357 12.11 59.52 ;
      END
   END FE_OFN53780_n_52084

   PIN FE_OFN53782_n_52084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.226 59.357 10.254 59.52 ;
      END
   END FE_OFN53782_n_52084

   PIN FE_OFN53783_n_52084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.514 59.357 22.542 59.52 ;
      END
   END FE_OFN53783_n_52084

   PIN FE_OFN53822_n_40455
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.586 0.163 33.614 ;
      END
   END FE_OFN53822_n_40455

   PIN FE_OFN53850_n_52081
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.178 59.357 16.206 59.52 ;
      END
   END FE_OFN53850_n_52081

   PIN FE_OFN53963_n_40967
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.834 0.163 30.862 ;
      END
   END FE_OFN53963_n_40967

   PIN FE_OFN53973_n_52082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.378 59.357 27.406 59.52 ;
      END
   END FE_OFN53973_n_52082

   PIN FE_OFN54887_n_45508
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 58.034 51.648 58.062 ;
      END
   END FE_OFN54887_n_45508

   PIN FE_OFN55725_n_52027
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 50.93 51.648 50.958 ;
      END
   END FE_OFN55725_n_52027

   PIN FE_OFN55732_n_52083
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.746 59.357 21.774 59.52 ;
      END
   END FE_OFN55732_n_52083

   PIN FE_OFN55733_n_52083
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.618 59.357 5.646 59.52 ;
      END
   END FE_OFN55733_n_52083

   PIN FE_OFN55736_n_52083
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.146 59.357 12.174 59.52 ;
      END
   END FE_OFN55736_n_52083

   PIN FE_OFN55761_n_52081
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.394 59.357 33.422 59.52 ;
      END
   END FE_OFN55761_n_52081

   PIN FE_OFN55822_n_52026
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.018 59.357 12.046 59.52 ;
      END
   END FE_OFN55822_n_52026

   PIN FE_OFN55823_n_52026
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.242 59.357 16.27 59.52 ;
      END
   END FE_OFN55823_n_52026

   PIN FE_OFN65159_n_57599
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 47.602 0.163 47.63 ;
      END
   END FE_OFN65159_n_57599

   PIN FE_OFN65264_n_40386
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.538 59.357 7.566 59.52 ;
      END
   END FE_OFN65264_n_40386

   PIN FE_OFN66190_n_40803
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 22.194 51.648 22.222 ;
      END
   END FE_OFN66190_n_40803

   PIN FE_OFN66462_n_41242
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.202 0.163 25.23 ;
      END
   END FE_OFN66462_n_41242

   PIN FE_OFN68662_n_41001
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.306 0.163 16.334 ;
      END
   END FE_OFN68662_n_41001

   PIN FE_OFN69662_n_40499
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.514 0.163 22.542 ;
      END
   END FE_OFN69662_n_40499

   PIN FE_OFN72075_n_35884
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.314 59.357 11.342 59.52 ;
      END
   END FE_OFN72075_n_35884

   PIN FE_OFN7415_n_57598
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.41 0.163 39.438 ;
      END
   END FE_OFN7415_n_57598

   PIN FE_OFN79894_n_53976
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.978 59.357 13.006 59.52 ;
      END
   END FE_OFN79894_n_53976

   PIN FE_OFN80051_n_54052
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 50.994 0.163 51.022 ;
      END
   END FE_OFN80051_n_54052

   PIN FE_OFN80076_n_57600
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.05 0.163 48.078 ;
      END
   END FE_OFN80076_n_57600

   PIN FE_OFN80128_n_40881
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.154 0.163 39.182 ;
      END
   END FE_OFN80128_n_40881

   PIN FE_OFN81050_n_40677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.21 0.163 20.238 ;
      END
   END FE_OFN81050_n_40677

   PIN FE_OFN82374_n_40595
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.162 0.163 2.19 ;
      END
   END FE_OFN82374_n_40595

   PIN FE_OFN89560_n_40600
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.186 0.163 43.214 ;
      END
   END FE_OFN89560_n_40600

   PIN FE_OFN89563_n_40669
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 33.65 0.163 33.678 ;
      END
   END FE_OFN89563_n_40669

   PIN FE_OFN89691_n_40666
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.85 0.163 36.878 ;
      END
   END FE_OFN89691_n_40666

   PIN FE_OFN89714_n_40740
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.514 0.163 30.542 ;
      END
   END FE_OFN89714_n_40740

   PIN FE_OFN89774_n_40818
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 38.642 0.163 38.67 ;
      END
   END FE_OFN89774_n_40818

   PIN FE_OFN89904_n_41210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.858 0.163 47.886 ;
      END
   END FE_OFN89904_n_41210

   PIN FE_OFN89935_n_40583
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.418 0.163 10.446 ;
      END
   END FE_OFN89935_n_40583

   PIN FE_OFN89944_n_40368
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END FE_OFN89944_n_40368

   PIN FE_OFN89967_n_40639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.794 0.163 47.822 ;
      END
   END FE_OFN89967_n_40639

   PIN FE_OFN89998_n_40672
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.818 59.357 24.846 59.52 ;
      END
   END FE_OFN89998_n_40672

   PIN FE_OFN90003_n_41246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.642 0.163 6.67 ;
      END
   END FE_OFN90003_n_41246

   PIN FE_OFN90026_n_40748
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.562 0.163 24.59 ;
      END
   END FE_OFN90026_n_40748

   PIN FE_OFN90039_n_40717
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.898 0.163 6.926 ;
      END
   END FE_OFN90039_n_40717

   PIN FE_OFN90040_n_40372
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.146 0.163 20.174 ;
      END
   END FE_OFN90040_n_40372

   PIN FE_OFN90041_n_40381
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.698 59.357 3.726 59.52 ;
      END
   END FE_OFN90041_n_40381

   PIN FE_OFN90067_n_40724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.042 0.163 45.07 ;
      END
   END FE_OFN90067_n_40724

   PIN FE_OFN90075_n_40436
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.986 59.357 16.014 59.52 ;
      END
   END FE_OFN90075_n_40436

   PIN FE_OFN90079_n_40674
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.882 59.357 16.91 59.52 ;
      END
   END FE_OFN90079_n_40674

   PIN FE_OFN90099_FE_OCPN63313_n_40689
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.25 0.163 11.278 ;
      END
   END FE_OFN90099_FE_OCPN63313_n_40689

   PIN FE_OFN92681_n_40584
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.018 0.163 20.046 ;
      END
   END FE_OFN92681_n_40584

   PIN FE_OFN92683_n_40586
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.61 0.163 42.638 ;
      END
   END FE_OFN92683_n_40586

   PIN FE_OFN92826_n_40562
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.762 0.163 27.79 ;
      END
   END FE_OFN92826_n_40562

   PIN FE_OFN92897_n_40742
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 43.122 0.163 43.15 ;
      END
   END FE_OFN92897_n_40742

   PIN FE_OFN93006_n_40725
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.09 0.163 7.118 ;
      END
   END FE_OFN93006_n_40725

   PIN FE_OFN93027_n_40885
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.33 0.163 25.358 ;
      END
   END FE_OFN93027_n_40885

   PIN FE_OFN93041_n_40615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.546 0.163 42.574 ;
      END
   END FE_OFN93041_n_40615

   PIN FE_OFN93057_n_40326
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.226 0.163 42.254 ;
      END
   END FE_OFN93057_n_40326

   PIN FE_OFN93058_n_40380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.602 0.163 15.63 ;
      END
   END FE_OFN93058_n_40380

   PIN FE_OFN93060_n_40468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.242 0.163 48.27 ;
      END
   END FE_OFN93060_n_40468

   PIN FE_OFN93171_n_40656
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 19.25 0.163 19.278 ;
      END
   END FE_OFN93171_n_40656

   PIN FE_OFN93173_n_41200
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.77 0.163 38.798 ;
      END
   END FE_OFN93173_n_41200

   PIN FE_OFN93186_n_40422
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.522 0.163 33.55 ;
      END
   END FE_OFN93186_n_40422

   PIN FE_OFN93289_n_40441
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.082 0.163 52.11 ;
      END
   END FE_OFN93289_n_40441

   PIN FE_OFN93291_n_40578
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.266 0.163 25.294 ;
      END
   END FE_OFN93291_n_40578

   PIN FE_OFN93292_n_40587
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.426 0.163 13.454 ;
      END
   END FE_OFN93292_n_40587

   PIN FE_OFN93294_n_40680
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.81 0.163 13.838 ;
      END
   END FE_OFN93294_n_40680

   PIN FE_OFN93352_n_40623
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 45.49 0.163 45.518 ;
      END
   END FE_OFN93352_n_40623

   PIN FE_OFN93353_n_40382
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.546 0.163 2.574 ;
      END
   END FE_OFN93353_n_40382

   PIN FE_OFN94636_n_40702
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.162 0.163 42.19 ;
      END
   END FE_OFN94636_n_40702

   PIN FE_OFN94776_n_40849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.698 0.163 11.726 ;
      END
   END FE_OFN94776_n_40849

   PIN FE_OFN94918_n_40413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.274 0.163 36.302 ;
      END
   END FE_OFN94918_n_40413

   PIN FE_OFN95014_n_41213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.09 0.163 39.118 ;
      END
   END FE_OFN95014_n_41213

   PIN FE_OFN95068_n_40835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.954 0.163 19.982 ;
      END
   END FE_OFN95068_n_40835

   PIN FE_OFN95079_n_40444
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.13 0.163 22.158 ;
      END
   END FE_OFN95079_n_40444

   PIN FE_OFN95120_n_40529
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.802 0.163 50.83 ;
      END
   END FE_OFN95120_n_40529

   PIN FE_OFN95165_n_40353
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 27.954 51.648 27.982 ;
      END
   END FE_OFN95165_n_40353

   PIN FE_OFN95201_n_40714
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.098 0.163 42.126 ;
      END
   END FE_OFN95201_n_40714

   PIN FE_OFN96060_FE_OCPN59260_n_40732
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.354 0.163 10.382 ;
      END
   END FE_OFN96060_FE_OCPN59260_n_40732

   PIN FE_OFN96766_FE_OCPN60886_n_40646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.066 0.163 22.094 ;
      END
   END FE_OFN96766_FE_OCPN60886_n_40646

   PIN FE_OFN96958_n_40592
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.73 0.163 47.758 ;
      END
   END FE_OFN96958_n_40592

   PIN FE_OFN97291_n_40798
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.57 0.163 27.598 ;
      END
   END FE_OFN97291_n_40798

   PIN FE_OFN97312_n_40440
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.002 0.163 22.03 ;
      END
   END FE_OFN97312_n_40440

   PIN FE_OFN97388_n_40734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.834 0.163 6.862 ;
      END
   END FE_OFN97388_n_40734

   PIN FE_OFN97595_FE_OCPN61185_n_40442
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.45 0.163 22.478 ;
      END
   END FE_OFN97595_FE_OCPN61185_n_40442

   PIN FE_RN_2180_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.25 59.357 35.278 59.52 ;
      END
   END FE_RN_2180_0

   PIN n_40316
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.698 0.163 27.726 ;
      END
   END n_40316

   PIN n_40337
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.706 0.163 38.734 ;
      END
   END n_40337

   PIN n_40354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.122 0.163 43.15 ;
      END
   END n_40354

   PIN n_40363
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.906 59.357 1.934 59.52 ;
      END
   END n_40363

   PIN n_40393
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.458 0.163 33.486 ;
      END
   END n_40393

   PIN n_40397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.77 0.163 6.798 ;
      END
   END n_40397

   PIN n_40404
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.034 0.163 42.062 ;
      END
   END n_40404

   PIN n_40409
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.97 0.163 41.998 ;
      END
   END n_40409

   PIN n_40414
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 42.29 0.163 42.318 ;
      END
   END n_40414

   PIN n_40418
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.178 0.163 48.206 ;
      END
   END n_40418

   PIN n_40423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.114 0.163 48.142 ;
      END
   END n_40423

   PIN n_40449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.57 0.163 11.598 ;
      END
   END n_40449

   PIN n_40460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.938 0.163 21.966 ;
      END
   END n_40460

   PIN n_40505
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.21 0.163 36.238 ;
      END
   END n_40505

   PIN n_40516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.362 59.357 5.39 59.52 ;
      END
   END n_40516

   PIN n_40526
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 43.25 0.163 43.278 ;
      END
   END n_40526

   PIN n_40556
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.514 59.357 30.542 59.52 ;
      END
   END n_40556

   PIN n_40579
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.506 0.163 11.534 ;
      END
   END n_40579

   PIN n_40593
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.026 0.163 39.054 ;
      END
   END n_40593

   PIN n_40598
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.642 0.163 38.67 ;
      END
   END n_40598

   PIN n_40616
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.666 0.163 47.694 ;
      END
   END n_40616

   PIN n_40637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.49 0.163 45.518 ;
      END
   END n_40637

   PIN n_40666
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.786 0.163 36.814 ;
      END
   END n_40666

   PIN n_40685
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.978 0.163 37.006 ;
      END
   END n_40685

   PIN n_40690
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 52.722 0.163 52.75 ;
      END
   END n_40690

   PIN n_40701
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.45 59.357 22.478 59.52 ;
      END
   END n_40701

   PIN n_40706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 36.53 0.163 36.558 ;
      END
   END n_40706

   PIN n_40710
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.906 0.163 41.934 ;
      END
   END n_40710

   PIN n_40720
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 45.426 0.163 45.454 ;
      END
   END n_40720

   PIN n_40729
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.002 59.357 6.03 59.52 ;
      END
   END n_40729

   PIN n_40741
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.506 59.357 27.534 59.52 ;
      END
   END n_40741

   PIN n_40743
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.394 0.163 33.422 ;
      END
   END n_40743

   PIN n_40745
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.226 0.163 34.254 ;
      END
   END n_40745

   PIN n_40765
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.146 0.163 36.174 ;
      END
   END n_40765

   PIN n_40768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 42.226 0.163 42.254 ;
      END
   END n_40768

   PIN n_40770
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.13 0.163 38.158 ;
      END
   END n_40770

   PIN n_40777
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.842 59.357 1.87 59.52 ;
      END
   END n_40777

   PIN n_40783
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.77 59.357 22.798 59.52 ;
      END
   END n_40783

   PIN n_41024
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.05 0.163 48.078 ;
      END
   END n_41024

   PIN n_41051
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.978 0.163 45.006 ;
      END
   END n_41051

   PIN n_41057
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 47.986 51.648 48.014 ;
      END
   END n_41057

   PIN n_41085
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.482 0.163 2.51 ;
      END
   END n_41085

   PIN n_41094
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.202 0.163 25.23 ;
      END
   END n_41094

   PIN n_41111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.45 0.163 30.478 ;
      END
   END n_41111

   PIN n_41129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.474 59.357 39.502 59.52 ;
      END
   END n_41129

   PIN n_41136
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 39.346 0.163 39.374 ;
      END
   END n_41136

   PIN n_41188
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.914 0.163 44.942 ;
      END
   END n_41188

   PIN n_41231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.946 0.163 24.974 ;
      END
   END n_41231

   PIN n_42980
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 51.485 39.41 51.648 39.438 ;
      END
   END n_42980

   PIN n_42981
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.97 59.357 41.998 59.52 ;
      END
   END n_42981

   PIN n_42983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.906 59.357 41.934 59.52 ;
      END
   END n_42983

   PIN n_45340
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.874 59.357 21.902 59.52 ;
      END
   END n_45340

   PIN n_45516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.85 59.357 44.878 59.52 ;
      END
   END n_45516

   PIN n_51367
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.69 59.357 48.718 59.52 ;
      END
   END n_51367

   PIN n_51369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.498 59.357 48.526 59.52 ;
      END
   END n_51369

   PIN n_53993
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.746 0.163 13.774 ;
      END
   END n_53993

   PIN n_54048
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.842 0.163 41.87 ;
      END
   END n_54048

   PIN n_54049
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.778 59.357 1.806 59.52 ;
      END
   END n_54049

   PIN n_54050
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.866 59.357 18.894 59.52 ;
      END
   END n_54050

   PIN n_54051
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.082 0.163 28.11 ;
      END
   END n_54051

   PIN n_54054
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.162 0.163 34.19 ;
      END
   END n_54054

   PIN n_54088
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.714 59.357 1.742 59.52 ;
      END
   END n_54088

   PIN n_54101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.85 0.163 44.878 ;
      END
   END n_54101

   PIN n_54219
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.594 59.357 4.622 59.52 ;
      END
   END n_54219

   PIN n_54222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.754 0.163 56.782 ;
      END
   END n_54222

   PIN n_56439
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 42.162 0.163 42.19 ;
      END
   END n_56439

   PIN n_57586
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.874 0.163 21.902 ;
      END
   END n_57586

   PIN n_58039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.058 59.357 19.086 59.52 ;
      END
   END n_58039

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 51.648 59.52 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 51.648 59.52 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 51.648 59.52 ;
      LAYER V1 ;
         RECT 0.0 0.0 51.648 59.52 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 51.648 59.52 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 51.648 59.52 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 51.648 59.52 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 51.648 59.52 ;
      LAYER M1 ;
         RECT 0.0 0.0 51.648 59.52 ;
   END
END h6_mgc_edit_dist_a

MACRO h3_mgc_edit_dist_a
   CLASS BLOCK ;
   FOREIGN h3 ;
   ORIGIN 0 0 ;
   SIZE 57.664 BY 64.64 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN56827_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.594 64.477 36.622 64.64 ;
      END
   END FE_OCPN56827_n_23035

   PIN FE_OCPN57195_FE_OFN46384_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.106 0.163 61.134 ;
      END
   END FE_OCPN57195_FE_OFN46384_n_23035

   PIN FE_OCPN57332_FE_OFN48190_n_22999
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 44.146 57.664 44.174 ;
      END
   END FE_OCPN57332_FE_OFN48190_n_22999

   PIN FE_OCPN58002_FE_OFN46384_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.17 0.163 61.198 ;
      END
   END FE_OCPN58002_FE_OFN46384_n_23035

   PIN FE_OCPN58799_FE_OFN41801_n_23039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.114 0.163 24.142 ;
      END
   END FE_OCPN58799_FE_OFN41801_n_23039

   PIN FE_OCPN59420_FE_OFN47458_n_22985
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.602 0.163 47.63 ;
      END
   END FE_OCPN59420_FE_OFN47458_n_22985

   PIN FE_OCPN59424_FE_OFN47458_n_22985
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 48.882 57.664 48.91 ;
      END
   END FE_OCPN59424_FE_OFN47458_n_22985

   PIN FE_OCPN59425_FE_OFN47458_n_22985
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.882 0.163 48.91 ;
      END
   END FE_OCPN59425_FE_OFN47458_n_22985

   PIN FE_OCPN59960_FE_OFN48190_n_22999
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 29.106 57.664 29.134 ;
      END
   END FE_OCPN59960_FE_OFN48190_n_22999

   PIN FE_OCPN60172_FE_OFN47326_n_67216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.81 0.163 29.838 ;
      END
   END FE_OCPN60172_FE_OFN47326_n_67216

   PIN FE_OCPN60404_FE_OFN48179_n_22997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 20.978 57.664 21.006 ;
      END
   END FE_OCPN60404_FE_OFN48179_n_22997

   PIN FE_OCPN61220_n_24492
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 26.994 57.664 27.022 ;
      END
   END FE_OCPN61220_n_24492

   PIN FE_OCPN61492_FE_OFN48190_n_22999
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.306 64.477 40.334 64.64 ;
      END
   END FE_OCPN61492_FE_OFN48190_n_22999

   PIN FE_OCPN63674_n_23815
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 49.522 57.664 49.55 ;
      END
   END FE_OCPN63674_n_23815

   PIN FE_OCPN76133_FE_OFN41801_n_23039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.178 0.163 24.206 ;
      END
   END FE_OCPN76133_FE_OFN41801_n_23039

   PIN FE_OCPN76840_FE_OFN47632_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.874 0.163 29.902 ;
      END
   END FE_OCPN76840_FE_OFN47632_n_22865

   PIN FE_OCPN76842_FE_OFN47632_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.658 0.0 12.686 0.163 ;
      END
   END FE_OCPN76842_FE_OFN47632_n_22865

   PIN FE_OCPN77030_FE_OFN75657_n_22948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.674 0.163 58.702 ;
      END
   END FE_OCPN77030_FE_OFN75657_n_22948

   PIN FE_OCP_RBN77248_FE_OCPN57193_FE_OFN46384_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.226 0.0 34.254 0.163 ;
      END
   END FE_OCP_RBN77248_FE_OCPN57193_FE_OFN46384_n_23035

   PIN FE_OCP_RBN77364_FE_OCPN57515_FE_OFN47099_n_23039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.042 0.0 53.07 0.163 ;
      END
   END FE_OCP_RBN77364_FE_OCPN57515_FE_OFN47099_n_23039

   PIN FE_OFN13351_n_25338
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.306 0.0 16.334 0.163 ;
      END
   END FE_OFN13351_n_25338

   PIN FE_OFN13710_n_23652
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.354 0.163 18.382 ;
      END
   END FE_OFN13710_n_23652

   PIN FE_OFN13716_n_24566
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 9.586 57.664 9.614 ;
      END
   END FE_OFN13716_n_24566

   PIN FE_OFN29431_n_522
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.194 0.0 22.222 0.163 ;
      END
   END FE_OFN29431_n_522

   PIN FE_OFN33789_n_3396
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.65 0.0 41.678 0.163 ;
      END
   END FE_OFN33789_n_3396

   PIN FE_OFN34206_n_82
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.13 0.0 22.158 0.163 ;
      END
   END FE_OFN34206_n_82

   PIN FE_OFN34223_n_81
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 32.69 57.664 32.718 ;
      END
   END FE_OFN34223_n_81

   PIN FE_OFN34312_n_77
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END FE_OFN34312_n_77

   PIN FE_OFN34580_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 7.154 57.664 7.182 ;
      END
   END FE_OFN34580_n_223

   PIN FE_OFN34592_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 12.722 57.664 12.75 ;
      END
   END FE_OFN34592_n_223

   PIN FE_OFN34595_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 36.082 57.664 36.11 ;
      END
   END FE_OFN34595_n_223

   PIN FE_OFN34606_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 21.234 57.664 21.262 ;
      END
   END FE_OFN34606_n_223

   PIN FE_OFN41924_n_227
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.418 0.163 18.446 ;
      END
   END FE_OFN41924_n_227

   PIN FE_OFN41991_n_228
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 38.45 57.664 38.478 ;
      END
   END FE_OFN41991_n_228

   PIN FE_OFN42299_n_47
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 12.594 57.664 12.622 ;
      END
   END FE_OFN42299_n_47

   PIN FE_OFN42492_n_33
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 49.074 57.664 49.102 ;
      END
   END FE_OFN42492_n_33

   PIN FE_OFN42501_n_33
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.282 0.0 55.31 0.163 ;
      END
   END FE_OFN42501_n_33

   PIN FE_OFN42529_n_32
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 41.33 57.664 41.358 ;
      END
   END FE_OFN42529_n_32

   PIN FE_OFN42808_n_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 18.418 57.664 18.446 ;
      END
   END FE_OFN42808_n_10

   PIN FE_OFN42954_n_3289
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 4.082 57.664 4.11 ;
      END
   END FE_OFN42954_n_3289

   PIN FE_OFN42968_n_1990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 52.786 57.664 52.814 ;
      END
   END FE_OFN42968_n_1990

   PIN FE_OFN43882_n_67219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.906 0.163 41.934 ;
      END
   END FE_OFN43882_n_67219

   PIN FE_OFN43982_mux_g_ln477_q_1311_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.626 0.0 8.654 0.163 ;
      END
   END FE_OFN43982_mux_g_ln477_q_1311_

   PIN FE_OFN47020_n_67217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.202 0.0 25.23 0.163 ;
      END
   END FE_OFN47020_n_67217

   PIN FE_OFN47329_n_67216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.754 0.163 32.782 ;
      END
   END FE_OFN47329_n_67216

   PIN FE_OFN47630_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.962 0.163 46.99 ;
      END
   END FE_OFN47630_n_22865

   PIN FE_OFN47632_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 21.234 57.664 21.262 ;
      END
   END FE_OFN47632_n_22865

   PIN FE_OFN48892_n_24195
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 12.53 57.664 12.558 ;
      END
   END FE_OFN48892_n_24195

   PIN FE_OFN51049_n_23652
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 32.562 57.664 32.59 ;
      END
   END FE_OFN51049_n_23652

   PIN FE_OFN51274_n_25014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 35.57 57.664 35.598 ;
      END
   END FE_OFN51274_n_25014

   PIN FE_OFN51275_n_25016
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 35.634 57.664 35.662 ;
      END
   END FE_OFN51275_n_25016

   PIN FE_OFN51548_n_23656
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 44.402 57.664 44.43 ;
      END
   END FE_OFN51548_n_23656

   PIN FE_OFN51552_n_23702
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 44.21 57.664 44.238 ;
      END
   END FE_OFN51552_n_23702

   PIN FE_OFN51947_n_23990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 61.042 57.664 61.07 ;
      END
   END FE_OFN51947_n_23990

   PIN FE_OFN52123_n_23549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 48.882 57.664 48.91 ;
      END
   END FE_OFN52123_n_23549

   PIN FE_OFN53748_n_3398
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.898 0.0 30.926 0.163 ;
      END
   END FE_OFN53748_n_3398

   PIN FE_OFN53753_n_71
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.29 64.477 42.318 64.64 ;
      END
   END FE_OFN53753_n_71

   PIN FE_OFN53899_n_89
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.778 0.0 49.806 0.163 ;
      END
   END FE_OFN53899_n_89

   PIN FE_OFN54457_n_23864
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.37 0.0 16.398 0.163 ;
      END
   END FE_OFN54457_n_23864

   PIN FE_OFN54621_n_23573
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 35.634 57.664 35.662 ;
      END
   END FE_OFN54621_n_23573

   PIN FE_OFN54630_n_23981
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 44.21 57.664 44.238 ;
      END
   END FE_OFN54630_n_23981

   PIN FE_OFN54631_n_23986
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 44.274 57.664 44.302 ;
      END
   END FE_OFN54631_n_23986

   PIN FE_OFN54638_n_24584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 38.578 57.664 38.606 ;
      END
   END FE_OFN54638_n_24584

   PIN FE_OFN54639_n_24584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.058 0.163 27.086 ;
      END
   END FE_OFN54639_n_24584

   PIN FE_OFN54891_n_23983
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 32.754 57.664 32.782 ;
      END
   END FE_OFN54891_n_23983

   PIN FE_OFN56004_n_5228837_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.682 0.163 61.71 ;
      END
   END FE_OFN56004_n_5228837_bar

   PIN FE_OFN71792_eq_15722_64_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.114 0.0 48.142 0.163 ;
      END
   END FE_OFN71792_eq_15722_64_n_18

   PIN FE_OFN73040_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 12.786 57.664 12.814 ;
      END
   END FE_OFN73040_n_23035

   PIN FE_OFN73486_n_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.186 0.0 35.214 0.163 ;
      END
   END FE_OFN73486_n_11

   PIN FE_OFN73506_n_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 61.362 57.664 61.39 ;
      END
   END FE_OFN73506_n_10

   PIN FE_OFN73546_n_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.594 0.0 36.622 0.163 ;
      END
   END FE_OFN73546_n_30

   PIN FE_OFN73612_n_43
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 48.946 57.664 48.974 ;
      END
   END FE_OFN73612_n_43

   PIN FE_OFN73633_n_31
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 11.058 57.664 11.086 ;
      END
   END FE_OFN73633_n_31

   PIN FE_OFN73665_n_33
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.218 64.477 55.246 64.64 ;
      END
   END FE_OFN73665_n_33

   PIN FE_OFN73711_n_222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.394 0.0 9.422 0.163 ;
      END
   END FE_OFN73711_n_222

   PIN FE_OFN74312_n_61
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.074 0.0 25.102 0.163 ;
      END
   END FE_OFN74312_n_61

   PIN FE_OFN75677_n_22920
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.842 0.163 49.87 ;
      END
   END FE_OFN75677_n_22920

   PIN FE_OFN81211_n_24583
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.49 0.0 13.518 0.163 ;
      END
   END FE_OFN81211_n_24583

   PIN FE_OFN85501_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.77 0.0 22.798 0.163 ;
      END
   END FE_OFN85501_n_223

   PIN FE_OFN86522_n_518
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.834 0.163 6.862 ;
      END
   END FE_OFN86522_n_518

   PIN FE_OFN87976_FE_OCPN56158_FE_OFN47027_n_67213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 48.242 57.664 48.27 ;
      END
   END FE_OFN87976_FE_OCPN56158_FE_OFN47027_n_67213

   PIN FE_OFN88160_n_22979
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.37 0.163 48.398 ;
      END
   END FE_OFN88160_n_22979

   PIN FE_OFN88164_n_22979
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.946 0.163 48.974 ;
      END
   END FE_OFN88164_n_22979

   PIN FE_OFN89154_n_865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.474 64.477 7.502 64.64 ;
      END
   END FE_OFN89154_n_865

   PIN FE_OFN90772_FE_OCPN60312_FE_OFN47628_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.01 0.163 49.038 ;
      END
   END FE_OFN90772_FE_OCPN60312_FE_OFN47628_n_22865

   PIN FE_OFN90794_n_22919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.802 0.163 50.83 ;
      END
   END FE_OFN90794_n_22919

   PIN FE_OFN90904_n_67217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.658 0.163 12.686 ;
      END
   END FE_OFN90904_n_67217

   PIN FE_OFN90954_FE_RN_2244_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 49.01 57.664 49.038 ;
      END
   END FE_OFN90954_FE_RN_2244_0

   PIN FE_OFN91045_n_25028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 48.306 57.664 48.334 ;
      END
   END FE_OFN91045_n_25028

   PIN FE_OFN93717_n_67217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.466 0.0 12.494 0.163 ;
      END
   END FE_OFN93717_n_67217

   PIN FE_OFN93911_n_23836
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 44.082 57.664 44.11 ;
      END
   END FE_OFN93911_n_23836

   PIN FE_OFN94059_n_23989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 55.794 57.664 55.822 ;
      END
   END FE_OFN94059_n_23989

   PIN FE_OFN94140_n_879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.17 64.477 53.198 64.64 ;
      END
   END FE_OFN94140_n_879

   PIN FE_OFN94180_FE_OCPN77031_FE_OFN75657_n_22948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.474 0.163 55.502 ;
      END
   END FE_OFN94180_FE_OCPN77031_FE_OFN75657_n_22948

   PIN FE_OFN98114_n_50
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.418 0.0 42.446 0.163 ;
      END
   END FE_OFN98114_n_50

   PIN FE_OFN98267_n_71
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.674 64.477 10.702 64.64 ;
      END
   END FE_OFN98267_n_71

   PIN FE_RN_4736_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.994 0.0 51.022 0.163 ;
      END
   END FE_RN_4736_0

   PIN FE_RN_4810_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 26.866 57.664 26.894 ;
      END
   END FE_RN_4810_0

   PIN FE_RN_5927_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 15.602 57.664 15.63 ;
      END
   END FE_RN_5927_0

   PIN mux_g_ln477_q_1304_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.786 0.0 52.814 0.163 ;
      END
   END mux_g_ln477_q_1304_

   PIN mux_g_ln477_q_1307_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 35.698 57.664 35.726 ;
      END
   END mux_g_ln477_q_1307_

   PIN mux_g_ln477_q_1311_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 56.306 57.664 56.334 ;
      END
   END mux_g_ln477_q_1311_

   PIN mux_g_ln477_q_1347_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.922 0.163 15.95 ;
      END
   END mux_g_ln477_q_1347_

   PIN mux_g_ln477_q_1350_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.914 0.0 4.942 0.163 ;
      END
   END mux_g_ln477_q_1350_

   PIN mux_g_ln477_q_1355_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 1.906 0.0 1.934 0.163 ;
      END
   END mux_g_ln477_q_1355_

   PIN mux_g_ln477_q_1364_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.098 0.0 2.126 0.163 ;
      END
   END mux_g_ln477_q_1364_

   PIN mux_g_ln477_q_1366_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.586 0.0 33.614 0.163 ;
      END
   END mux_g_ln477_q_1366_

   PIN mux_g_ln477_q_1480_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.986 0.163 24.014 ;
      END
   END mux_g_ln477_q_1480_

   PIN mux_g_ln477_q_1484_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 44.338 57.664 44.366 ;
      END
   END mux_g_ln477_q_1484_

   PIN mux_g_ln477_q_1488_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.858 0.0 7.886 0.163 ;
      END
   END mux_g_ln477_q_1488_

   PIN mux_g_ln477_q_1496_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.026 0.163 47.054 ;
      END
   END mux_g_ln477_q_1496_

   PIN mux_g_ln477_q_1497_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.802 0.163 34.83 ;
      END
   END mux_g_ln477_q_1497_

   PIN mux_g_ln477_q_1500_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 29.17 57.664 29.198 ;
      END
   END mux_g_ln477_q_1500_

   PIN mux_g_ln477_q_1503_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.914 0.163 52.942 ;
      END
   END mux_g_ln477_q_1503_

   PIN mux_g_ln477_q_1534_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.202 64.477 25.23 64.64 ;
      END
   END mux_g_ln477_q_1534_

   PIN mux_g_ln477_q_578_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.834 0.0 54.862 0.163 ;
      END
   END mux_g_ln477_q_578_

   PIN mux_g_ln477_q_592_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.93 0.0 26.958 0.163 ;
      END
   END mux_g_ln477_q_592_

   PIN mux_g_ln477_q_593_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.434 0.0 16.462 0.163 ;
      END
   END mux_g_ln477_q_593_

   PIN mux_g_ln477_q_597_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.714 0.0 33.742 0.163 ;
      END
   END mux_g_ln477_q_597_

   PIN mux_g_ln477_q_601_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.778 0.0 33.806 0.163 ;
      END
   END mux_g_ln477_q_601_

   PIN mux_g_ln477_q_602_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.066 0.0 22.094 0.163 ;
      END
   END mux_g_ln477_q_602_

   PIN mux_g_ln477_q_604_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.858 0.0 31.886 0.163 ;
      END
   END mux_g_ln477_q_604_

   PIN n_2109
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.874 0.0 53.902 0.163 ;
      END
   END n_2109

   PIN n_2226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 24.178 57.664 24.206 ;
      END
   END n_2226

   PIN n_23565
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.97 0.163 49.998 ;
      END
   END n_23565

   PIN n_23712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 3.442 57.664 3.47 ;
      END
   END n_23712

   PIN n_23850
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 27.122 57.664 27.15 ;
      END
   END n_23850

   PIN n_23872
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 16.37 57.664 16.398 ;
      END
   END n_23872

   PIN n_23898
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 47.09 57.664 47.118 ;
      END
   END n_23898

   PIN n_23911
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 21.106 57.664 21.134 ;
      END
   END n_23911

   PIN n_24578
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 41.842 57.664 41.87 ;
      END
   END n_24578

   PIN n_24650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 22.514 57.664 22.542 ;
      END
   END n_24650

   PIN n_24655
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 12.466 57.664 12.494 ;
      END
   END n_24655

   PIN n_24658
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.89 0.0 27.918 0.163 ;
      END
   END n_24658

   PIN n_24848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 7.026 57.664 7.054 ;
      END
   END n_24848

   PIN n_25026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 48.37 57.664 48.398 ;
      END
   END n_25026

   PIN n_25030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.674 0.0 10.702 0.163 ;
      END
   END n_25030

   PIN n_25035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.354 64.477 42.382 64.64 ;
      END
   END n_25035

   PIN n_25044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.034 0.163 50.062 ;
      END
   END n_25044

   PIN n_25299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 29.682 57.664 29.71 ;
      END
   END n_25299

   PIN n_25309
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 32.882 57.664 32.91 ;
      END
   END n_25309

   PIN n_2712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 7.026 57.664 7.054 ;
      END
   END n_2712

   PIN n_2800
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.946 0.0 24.974 0.163 ;
      END
   END n_2800

   PIN n_2812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 2.866 57.664 2.894 ;
      END
   END n_2812

   PIN n_3110
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 21.042 57.664 21.07 ;
      END
   END n_3110

   PIN n_3283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 2.802 57.664 2.83 ;
      END
   END n_3283

   PIN n_3290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.874 0.0 53.902 0.163 ;
      END
   END n_3290

   PIN n_4733
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.818 0.163 32.846 ;
      END
   END n_4733

   PIN n_5562
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.042 0.0 13.07 0.163 ;
      END
   END n_5562

   PIN n_5563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.402 0.0 4.43 0.163 ;
      END
   END n_5563

   PIN n_5890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.906 0.163 9.934 ;
      END
   END n_5890

   PIN n_6316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.514 0.163 22.542 ;
      END
   END n_6316

   PIN n_6739
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.178 0.0 48.206 0.163 ;
      END
   END n_6739

   PIN FE_OCPN56158_FE_OFN47027_n_67213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 45.042 57.664 45.07 ;
      END
   END FE_OCPN56158_FE_OFN47027_n_67213

   PIN FE_OCPN56824_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 42.482 57.664 42.51 ;
      END
   END FE_OCPN56824_n_23035

   PIN FE_OCPN57568_FE_OFN47196_n_67214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.882 0.0 24.91 0.163 ;
      END
   END FE_OCPN57568_FE_OFN47196_n_67214

   PIN FE_OCPN58871_FE_OFN43374_n_22937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 29.81 57.664 29.838 ;
      END
   END FE_OCPN58871_FE_OFN43374_n_22937

   PIN FE_OCPN59418_FE_OFN47458_n_22985
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 7.09 57.664 7.118 ;
      END
   END FE_OCPN59418_FE_OFN47458_n_22985

   PIN FE_OCPN59878_FE_OFN47327_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 18.354 57.664 18.382 ;
      END
   END FE_OCPN59878_FE_OFN47327_n_67216

   PIN FE_OCPN59929_FE_OFN47456_n_22985
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 27.058 57.664 27.086 ;
      END
   END FE_OCPN59929_FE_OFN47456_n_22985

   PIN FE_OCPN59934_n_24570
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 15.282 57.664 15.31 ;
      END
   END FE_OCPN59934_n_24570

   PIN FE_OCPN60169_FE_OFN47326_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 6.834 57.664 6.862 ;
      END
   END FE_OCPN60169_FE_OFN47326_n_67216

   PIN FE_OCPN60170_FE_OFN47326_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 9.97 57.664 9.998 ;
      END
   END FE_OCPN60170_FE_OFN47326_n_67216

   PIN FE_OCPN60246_FE_OFN47005_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 18.546 57.664 18.574 ;
      END
   END FE_OCPN60246_FE_OFN47005_n_67217

   PIN FE_OCPN60333_FE_OFN41824_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 39.282 57.664 39.31 ;
      END
   END FE_OCPN60333_FE_OFN41824_n_23039

   PIN FE_OCPN60351_FE_OFN43508_n_22865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.29 0.0 42.318 0.163 ;
      END
   END FE_OCPN60351_FE_OFN43508_n_22865

   PIN FE_OCPN60402_FE_OFN48179_n_22997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 19.442 57.664 19.47 ;
      END
   END FE_OCPN60402_FE_OFN48179_n_22997

   PIN FE_OCPN61219_n_24492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.122 64.477 11.15 64.64 ;
      END
   END FE_OCPN61219_n_24492

   PIN FE_OCPN63510_FE_OFN41801_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 12.658 57.664 12.686 ;
      END
   END FE_OCPN63510_FE_OFN41801_n_23039

   PIN FE_OCPN77813_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 18.482 57.664 18.51 ;
      END
   END FE_OCPN77813_n_23035

   PIN FE_OCPN77821_FE_OFN47978_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.65 0.0 33.678 0.163 ;
      END
   END FE_OCPN77821_FE_OFN47978_n_23035

   PIN FE_OCPN77894_n_23972
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 54.066 57.664 54.094 ;
      END
   END FE_OCPN77894_n_23972

   PIN FE_OCPN78264_FE_OFN47649_n_22866
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.842 0.0 41.87 0.163 ;
      END
   END FE_OCPN78264_FE_OFN47649_n_22866

   PIN FE_OCPN95395_FE_OFN46375_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 21.17 57.664 21.198 ;
      END
   END FE_OCPN95395_FE_OFN46375_n_23035

   PIN FE_OCPN95638_FE_OFN48190_n_22999
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 16.306 57.664 16.334 ;
      END
   END FE_OCPN95638_FE_OFN48190_n_22999

   PIN FE_OCPUNCON99093_FE_OCP_RBN77363_FE_OCPN57515_FE_OFN47099_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.73 64.477 7.758 64.64 ;
      END
   END FE_OCPUNCON99093_FE_OCP_RBN77363_FE_OCPN57515_FE_OFN47099_n_23039

   PIN FE_OCP_RBN77173_FE_OFN46375_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.426 0.0 29.454 0.163 ;
      END
   END FE_OCP_RBN77173_FE_OFN46375_n_23035

   PIN FE_OFN13154_n_25272
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 22.45 57.664 22.478 ;
      END
   END FE_OFN13154_n_25272

   PIN FE_OFN13349_n_25338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 9.522 57.664 9.55 ;
      END
   END FE_OFN13349_n_25338

   PIN FE_OFN15344_n_24443
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 16.242 57.664 16.27 ;
      END
   END FE_OFN15344_n_24443

   PIN FE_OFN29701_n_518
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.81 0.0 21.838 0.163 ;
      END
   END FE_OFN29701_n_518

   PIN FE_OFN34029_n_89
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.866 64.477 42.894 64.64 ;
      END
   END FE_OFN34029_n_89

   PIN FE_OFN34082_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.314 0.0 19.342 0.163 ;
      END
   END FE_OFN34082_n_87

   PIN FE_OFN34202_n_82
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 36.21 57.664 36.238 ;
      END
   END FE_OFN34202_n_82

   PIN FE_OFN34291_n_78
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 54.13 57.664 54.158 ;
      END
   END FE_OFN34291_n_78

   PIN FE_OFN34467_n_59
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.386 0.0 46.414 0.163 ;
      END
   END FE_OFN34467_n_59

   PIN FE_OFN34549_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 29.234 57.664 29.262 ;
      END
   END FE_OFN34549_n_223

   PIN FE_OFN34560_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.01 0.0 25.038 0.163 ;
      END
   END FE_OFN34560_n_223

   PIN FE_OFN35094_n_5228270_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.626 64.477 40.654 64.64 ;
      END
   END FE_OFN35094_n_5228270_bar

   PIN FE_OFN35482_eq_15722_64_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.154 64.477 55.182 64.64 ;
      END
   END FE_OFN35482_eq_15722_64_n_18

   PIN FE_OFN42005_n_231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.226 64.477 18.254 64.64 ;
      END
   END FE_OFN42005_n_231

   PIN FE_OFN42081_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.498 0.0 32.526 0.163 ;
      END
   END FE_OFN42081_n_222

   PIN FE_OFN42082_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.426 0.0 13.454 0.163 ;
      END
   END FE_OFN42082_n_222

   PIN FE_OFN42113_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.498 64.477 48.526 64.64 ;
      END
   END FE_OFN42113_n_222

   PIN FE_OFN42143_n_57
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.194 64.477 22.222 64.64 ;
      END
   END FE_OFN42143_n_57

   PIN FE_OFN42297_n_47
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 35.506 57.664 35.534 ;
      END
   END FE_OFN42297_n_47

   PIN FE_OFN42346_n_45
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 44.274 57.664 44.302 ;
      END
   END FE_OFN42346_n_45

   PIN FE_OFN42388_n_43
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.378 64.477 19.406 64.64 ;
      END
   END FE_OFN42388_n_43

   PIN FE_OFN42435_n_41
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.874 64.477 45.902 64.64 ;
      END
   END FE_OFN42435_n_41

   PIN FE_OFN42544_n_31
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.402 64.477 44.43 64.64 ;
      END
   END FE_OFN42544_n_31

   PIN FE_OFN42570_n_30
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.042 64.477 37.07 64.64 ;
      END
   END FE_OFN42570_n_30

   PIN FE_OFN42595_n_29
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.25 64.477 19.278 64.64 ;
      END
   END FE_OFN42595_n_29

   PIN FE_OFN42596_n_29
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.314 64.477 19.342 64.64 ;
      END
   END FE_OFN42596_n_29

   PIN FE_OFN42629_n_20
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 48.242 57.664 48.27 ;
      END
   END FE_OFN42629_n_20

   PIN FE_OFN42789_n_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 29.042 57.664 29.07 ;
      END
   END FE_OFN42789_n_11

   PIN FE_OFN42953_n_3289
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.594 0.163 12.622 ;
      END
   END FE_OFN42953_n_3289

   PIN FE_OFN43845_n_67218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.45 0.0 14.478 0.082 ;
      END
   END FE_OFN43845_n_67218

   PIN FE_OFN43847_n_67218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.786 0.0 4.814 0.082 ;
      END
   END FE_OFN43847_n_67218

   PIN FE_OFN46995_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 24.114 57.664 24.142 ;
      END
   END FE_OFN46995_n_67217

   PIN FE_OFN46996_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 22.578 57.664 22.606 ;
      END
   END FE_OFN46996_n_67217

   PIN FE_OFN47017_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.114 0.0 48.142 0.163 ;
      END
   END FE_OFN47017_n_67217

   PIN FE_OFN47019_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.002 0.0 38.03 0.163 ;
      END
   END FE_OFN47019_n_67217

   PIN FE_OFN47328_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 22.002 57.664 22.03 ;
      END
   END FE_OFN47328_n_67216

   PIN FE_OFN47628_n_22865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 48.434 57.664 48.462 ;
      END
   END FE_OFN47628_n_22865

   PIN FE_OFN47808_n_22977
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.842 0.0 17.87 0.163 ;
      END
   END FE_OFN47808_n_22977

   PIN FE_OFN47977_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.65 0.0 33.678 0.163 ;
      END
   END FE_OFN47977_n_23035

   PIN FE_OFN48729_n_865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.738 0.163 58.766 ;
      END
   END FE_OFN48729_n_865

   PIN FE_OFN48776_n_879
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.954 0.0 27.982 0.163 ;
      END
   END FE_OFN48776_n_879

   PIN FE_OFN50050_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.69 0.0 16.718 0.082 ;
      END
   END FE_OFN50050_n_71

   PIN FE_OFN51564_n_23989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.306 0.163 48.334 ;
      END
   END FE_OFN51564_n_23989

   PIN FE_OFN51946_n_23990
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.042 0.163 61.07 ;
      END
   END FE_OFN51946_n_23990

   PIN FE_OFN53694_n_91
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.45 0.163 22.478 ;
      END
   END FE_OFN53694_n_91

   PIN FE_OFN53750_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.402 64.477 28.43 64.64 ;
      END
   END FE_OFN53750_n_71

   PIN FE_OFN53910_n_77
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 9.906 57.664 9.934 ;
      END
   END FE_OFN53910_n_77

   PIN FE_OFN53911_n_77
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.514 0.0 54.542 0.163 ;
      END
   END FE_OFN53911_n_77

   PIN FE_OFN72259_n_3398
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.946 64.477 48.974 64.64 ;
      END
   END FE_OFN72259_n_3398

   PIN FE_OFN73407_n_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 36.146 57.664 36.174 ;
      END
   END FE_OFN73407_n_14

   PIN FE_OFN73437_n_40
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.93 0.163 26.958 ;
      END
   END FE_OFN73437_n_40

   PIN FE_OFN73503_n_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.898 64.477 54.926 64.64 ;
      END
   END FE_OFN73503_n_10

   PIN FE_OFN73527_n_42
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 32.818 57.664 32.846 ;
      END
   END FE_OFN73527_n_42

   PIN FE_OFN73542_n_30
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 23.986 57.664 24.014 ;
      END
   END FE_OFN73542_n_30

   PIN FE_OFN73592_n_44
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.53 64.477 36.558 64.64 ;
      END
   END FE_OFN73592_n_44

   PIN FE_OFN73597_n_44
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 41.906 57.664 41.934 ;
      END
   END FE_OFN73597_n_44

   PIN FE_OFN73753_n_227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 6.962 57.664 6.99 ;
      END
   END FE_OFN73753_n_227

   PIN FE_OFN74310_n_61
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 47.026 57.664 47.054 ;
      END
   END FE_OFN74310_n_61

   PIN FE_OFN74425_n_81
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 18.354 57.664 18.382 ;
      END
   END FE_OFN74425_n_81

   PIN FE_OFN74585_n_79
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 29.426 57.664 29.454 ;
      END
   END FE_OFN74585_n_79

   PIN FE_OFN74729_n_522
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.05 0.163 24.078 ;
      END
   END FE_OFN74729_n_522

   PIN FE_OFN74760_n_528
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.234 0.0 13.262 0.163 ;
      END
   END FE_OFN74760_n_528

   PIN FE_OFN75614_n_67219
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.394 64.477 33.422 64.64 ;
      END
   END FE_OFN75614_n_67219

   PIN FE_OFN79568_n_24853
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 9.842 57.664 9.87 ;
      END
   END FE_OFN79568_n_24853

   PIN FE_OFN81210_n_24583
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 23.282 57.664 23.31 ;
      END
   END FE_OFN81210_n_24583

   PIN FE_OFN85037_n_16
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.306 64.477 32.334 64.64 ;
      END
   END FE_OFN85037_n_16

   PIN FE_OFN85123_n_33
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.018 0.0 28.046 0.163 ;
      END
   END FE_OFN85123_n_33

   PIN FE_OFN85133_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 32.626 57.664 32.654 ;
      END
   END FE_OFN85133_n_222

   PIN FE_OFN85161_n_228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.338 64.477 52.366 64.64 ;
      END
   END FE_OFN85161_n_228

   PIN FE_OFN88159_n_22979
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.074 64.477 25.102 64.64 ;
      END
   END FE_OFN88159_n_22979

   PIN FE_OFN88474_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 18.29 57.664 18.318 ;
      END
   END FE_OFN88474_n_23035

   PIN FE_OFN90605_n_22920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 52.914 57.664 52.942 ;
      END
   END FE_OFN90605_n_22920

   PIN FE_OFN90793_n_22919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 50.802 57.664 50.83 ;
      END
   END FE_OFN90793_n_22919

   PIN FE_OFN91248_n_22948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.501 52.914 57.664 52.942 ;
      END
   END FE_OFN91248_n_22948

   PIN FE_OFN91275_n_24566
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 16.818 57.664 16.846 ;
      END
   END FE_OFN91275_n_24566

   PIN FE_OFN91539_n_24449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 38.514 57.664 38.542 ;
      END
   END FE_OFN91539_n_24449

   PIN FE_OFN93720_n_22938
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.842 0.163 41.87 ;
      END
   END FE_OFN93720_n_22938

   PIN FE_OFN94058_n_23983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.794 0.0 7.822 0.163 ;
      END
   END FE_OFN94058_n_23983

   PIN FE_OFN98113_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.042 0.163 29.07 ;
      END
   END FE_OFN98113_n_50

   PIN FE_OFN98889_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.17 0.0 45.198 0.163 ;
      END
   END FE_OFN98889_n_67217

   PIN FE_RN_2244_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 18.226 57.664 18.254 ;
      END
   END FE_RN_2244_0

   PIN FE_RN_4805_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.034 0.0 2.062 0.163 ;
      END
   END FE_RN_4805_0

   PIN a_in_203_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 41.394 0.163 41.422 ;
      END
   END a_in_203_0

   PIN a_in_208_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.066 0.163 30.094 ;
      END
   END a_in_208_0

   PIN a_in_208_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.538 0.163 15.566 ;
      END
   END a_in_208_3

   PIN a_in_209_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.458 0.163 41.486 ;
      END
   END a_in_209_2

   PIN a_in_20_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.378 0.0 19.406 0.163 ;
      END
   END a_in_20_0

   PIN a_in_20_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 29.874 0.163 29.902 ;
      END
   END a_in_20_1

   PIN a_in_20_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.018 0.163 4.046 ;
      END
   END a_in_20_2

   PIN a_in_20_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.298 0.163 21.326 ;
      END
   END a_in_20_3

   PIN a_in_210_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 41.33 0.163 41.358 ;
      END
   END a_in_210_2

   PIN a_in_210_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.394 0.163 41.422 ;
      END
   END a_in_210_3

   PIN a_in_213_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 61.554 0.163 61.582 ;
      END
   END a_in_213_0

   PIN a_in_22_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.474 0.163 15.502 ;
      END
   END a_in_22_0

   PIN a_in_22_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.986 0.0 40.014 0.163 ;
      END
   END a_in_22_1

   PIN a_in_23_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.354 0.0 42.382 0.163 ;
      END
   END a_in_23_0

   PIN a_in_242_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 47.346 0.163 47.374 ;
      END
   END a_in_242_2

   PIN a_in_243_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.282 0.163 47.31 ;
      END
   END a_in_243_2

   PIN a_in_246_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 35.634 0.163 35.662 ;
      END
   END a_in_246_1

   PIN a_in_247_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.746 0.163 29.774 ;
      END
   END a_in_247_1

   PIN a_in_251_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.73 0.163 55.758 ;
      END
   END a_in_251_2

   PIN a_in_253_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.474 0.0 39.502 0.163 ;
      END
   END a_in_253_1

   PIN a_in_253_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.266 0.163 41.294 ;
      END
   END a_in_253_2

   PIN a_in_255_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.298 0.163 61.326 ;
      END
   END a_in_255_2

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.714 0.082 9.742 ;
      END
   END ispd_clk

   PIN memread_edit_dist_g2_ln254_unr113_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.674 0.0 10.702 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr113_q_6_

   PIN memread_edit_dist_g2_ln254_unr48_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.834 0.0 30.862 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr48_q_0_

   PIN memread_edit_dist_g2_ln254_unr48_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.218 0.0 55.246 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr48_q_4_

   PIN memread_edit_dist_g2_ln254_unr49_q_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.954 0.0 27.982 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_10_

   PIN memread_edit_dist_g2_ln254_unr49_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.506 0.0 35.534 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_1_

   PIN memread_edit_dist_g2_ln254_unr49_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.338 0.0 52.366 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_2_

   PIN memread_edit_dist_g2_ln254_unr49_q_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.922 0.0 23.95 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_3_

   PIN memread_edit_dist_g2_ln254_unr49_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.666 0.0 7.694 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_6_

   PIN memread_edit_dist_g2_ln254_unr49_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.73 0.0 7.758 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_7_

   PIN memread_edit_dist_g2_ln254_unr49_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.418 0.0 10.446 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_8_

   PIN mux_g_ln477_q_1324_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.178 0.0 48.206 0.163 ;
      END
   END mux_g_ln477_q_1324_

   PIN mux_g_ln477_q_1344_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.538 0.0 15.566 0.163 ;
      END
   END mux_g_ln477_q_1344_

   PIN mux_g_ln477_q_1354_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.994 0.163 27.022 ;
      END
   END mux_g_ln477_q_1354_

   PIN mux_g_ln477_q_1481_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 35.378 57.664 35.406 ;
      END
   END mux_g_ln477_q_1481_

   PIN mux_g_ln477_q_1482_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.242 0.163 48.27 ;
      END
   END mux_g_ln477_q_1482_

   PIN mux_g_ln477_q_1486_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.338 0.163 44.366 ;
      END
   END mux_g_ln477_q_1486_

   PIN mux_g_ln477_q_1501_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.906 0.163 49.934 ;
      END
   END mux_g_ln477_q_1501_

   PIN mux_g_ln477_q_1518_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.162 64.477 2.19 64.64 ;
      END
   END mux_g_ln477_q_1518_

   PIN mux_g_ln477_q_1525_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.914 64.477 4.942 64.64 ;
      END
   END mux_g_ln477_q_1525_

   PIN mux_g_ln477_q_1526_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.61 0.0 10.638 0.163 ;
      END
   END mux_g_ln477_q_1526_

   PIN mux_g_ln477_q_600_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.85 0.0 20.878 0.163 ;
      END
   END mux_g_ln477_q_600_

   PIN n_1788
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.578 0.163 38.606 ;
      END
   END n_1788

   PIN n_1861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.138 0.0 25.166 0.163 ;
      END
   END n_1861

   PIN n_1990
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.426 0.0 45.454 0.163 ;
      END
   END n_1990

   PIN n_2013
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.354 0.0 50.382 0.163 ;
      END
   END n_2013

   PIN n_2044
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.834 0.0 30.862 0.163 ;
      END
   END n_2044

   PIN n_2050
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.514 0.163 38.542 ;
      END
   END n_2050

   PIN n_2070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.034 0.0 2.062 0.163 ;
      END
   END n_2070

   PIN n_2108
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.466 0.0 20.494 0.163 ;
      END
   END n_2108

   PIN n_2202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 6.898 57.664 6.926 ;
      END
   END n_2202

   PIN n_2260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.066 0.163 54.094 ;
      END
   END n_2260

   PIN n_23549
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.274 0.163 44.302 ;
      END
   END n_23549

   PIN n_23573
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.194 0.0 6.222 0.163 ;
      END
   END n_23573

   PIN n_23650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.97 0.163 9.998 ;
      END
   END n_23650

   PIN n_23702
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.482 0.163 42.51 ;
      END
   END n_23702

   PIN n_23746
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.578 0.163 22.606 ;
      END
   END n_23746

   PIN n_23815
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.85 0.163 52.878 ;
      END
   END n_23815

   PIN n_23843
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 26.994 57.664 27.022 ;
      END
   END n_23843

   PIN n_23864
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.578 0.0 14.606 0.163 ;
      END
   END n_23864

   PIN n_23901
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 54.002 57.664 54.03 ;
      END
   END n_23901

   PIN n_23981
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.634 0.163 35.662 ;
      END
   END n_23981

   PIN n_23986
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.202 0.163 41.23 ;
      END
   END n_23986

   PIN n_2402
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.498 0.0 16.526 0.163 ;
      END
   END n_2402

   PIN n_2412
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.53 0.0 36.558 0.163 ;
      END
   END n_2412

   PIN n_24195
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.226 0.0 42.254 0.163 ;
      END
   END n_24195

   PIN n_24445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 29.746 57.664 29.774 ;
      END
   END n_24445

   PIN n_24462
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 24.05 57.664 24.078 ;
      END
   END n_24462

   PIN n_24465
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 18.162 57.664 18.19 ;
      END
   END n_24465

   PIN n_2450
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 49.842 57.664 49.87 ;
      END
   END n_2450

   PIN n_24851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.706 0.0 30.734 0.163 ;
      END
   END n_24851

   PIN n_24855
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 26.93 57.664 26.958 ;
      END
   END n_24855

   PIN n_25014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.57 0.163 35.598 ;
      END
   END n_25014

   PIN n_25016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.45 0.163 38.478 ;
      END
   END n_25016

   PIN n_2513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.842 0.163 9.87 ;
      END
   END n_2513

   PIN n_25319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 35.442 57.664 35.47 ;
      END
   END n_25319

   PIN n_2593
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.77 0.0 30.798 0.163 ;
      END
   END n_2593

   PIN n_2628
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.33 0.0 9.358 0.163 ;
      END
   END n_2628

   PIN n_2642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.45 0.0 46.478 0.163 ;
      END
   END n_2642

   PIN n_2754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.898 0.163 6.926 ;
      END
   END n_2754

   PIN n_2809
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.77 0.163 22.798 ;
      END
   END n_2809

   PIN n_2826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.002 0.163 54.03 ;
      END
   END n_2826

   PIN n_2944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.506 0.163 35.534 ;
      END
   END n_2944

   PIN n_2986
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.442 0.163 3.47 ;
      END
   END n_2986

   PIN n_3111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.29 0.163 18.318 ;
      END
   END n_3111

   PIN n_3265
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.954 0.163 3.982 ;
      END
   END n_3265

   PIN n_3303
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.074 0.0 25.102 0.163 ;
      END
   END n_3303

   PIN n_48
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.442 0.163 35.47 ;
      END
   END n_48

   PIN n_5228837_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.562 64.477 8.59 64.64 ;
      END
   END n_5228837_bar

   PIN n_5347
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.602 0.163 15.63 ;
      END
   END n_5347

   PIN n_5409
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.058 64.477 43.086 64.64 ;
      END
   END n_5409

   PIN n_6457
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.501 52.85 57.664 52.878 ;
      END
   END n_6457

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 57.664 64.64 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 57.664 64.64 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 57.664 64.64 ;
      LAYER V1 ;
         RECT 0.0 0.0 57.664 64.64 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 57.664 64.64 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 57.664 64.64 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 57.664 64.64 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 57.664 64.64 ;
      LAYER M1 ;
         RECT 0.0 0.0 57.664 64.64 ;
   END
END h3_mgc_edit_dist_a

MACRO h2_mgc_edit_dist_a
   CLASS BLOCK ;
   FOREIGN h2 ;
   ORIGIN 0 0 ;
   SIZE 57.728 BY 37.12 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN61466_FE_OFN48299_n_31625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.565 10.354 57.728 10.382 ;
      END
   END FE_OCPN61466_FE_OFN48299_n_31625

   PIN FE_OCPN78682_n_32759
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.818 0.163 24.846 ;
      END
   END FE_OCPN78682_n_32759

   PIN FE_OCPN99272_FE_OFN46361_n_67216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.042 0.0 13.07 0.163 ;
      END
   END FE_OCPN99272_FE_OFN46361_n_67216

   PIN FE_OCPUNCON78515_ternarymux_ln49_0_unr82_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 13.17 57.728 13.198 ;
      END
   END FE_OCPUNCON78515_ternarymux_ln49_0_unr82_z_3_

   PIN FE_OFN30000_n_35944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 27.186 0.163 27.214 ;
      END
   END FE_OFN30000_n_35944

   PIN FE_OFN30327_n_36003
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.93 0.163 18.958 ;
      END
   END FE_OFN30327_n_36003

   PIN FE_OFN30401_n_35970
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.482 0.163 10.51 ;
      END
   END FE_OFN30401_n_35970

   PIN FE_OFN30534_n_36241
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.866 0.163 18.894 ;
      END
   END FE_OFN30534_n_36241

   PIN FE_OFN30638_n_36637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.834 0.163 22.862 ;
      END
   END FE_OFN30638_n_36637

   PIN FE_OFN35164_memwrite_edit_dist_g2_ln280_unr61_en_0__4469706
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.13 0.163 6.158 ;
      END
   END FE_OFN35164_memwrite_edit_dist_g2_ln280_unr61_en_0__4469706

   PIN FE_OFN42686_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 2.418 57.728 2.446 ;
      END
   END FE_OFN42686_n_15

   PIN FE_OFN42687_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.762 36.957 51.79 37.12 ;
      END
   END FE_OFN42687_n_15

   PIN FE_OFN42689_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.898 0.0 54.926 0.163 ;
      END
   END FE_OFN42689_n_15

   PIN FE_OFN42935_n_2966
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.794 0.0 47.822 0.163 ;
      END
   END FE_OFN42935_n_2966

   PIN FE_OFN46788_n_26948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.81 0.163 5.838 ;
      END
   END FE_OFN46788_n_26948

   PIN FE_OFN49891_n_93
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.77 0.0 54.798 0.163 ;
      END
   END FE_OFN49891_n_93

   PIN FE_OFN53694_n_91
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.226 0.163 2.254 ;
      END
   END FE_OFN53694_n_91

   PIN FE_OFN54144_ternarymux_ln49_0_unr61_z_10__4330982
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.882 0.163 24.91 ;
      END
   END FE_OFN54144_ternarymux_ln49_0_unr61_z_10__4330982

   PIN FE_OFN54360_memread_edit_dist_a_ln268_unr124_a_33__4330321
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 2.226 57.728 2.254 ;
      END
   END FE_OFN54360_memread_edit_dist_a_ln268_unr124_a_33__4330321

   PIN FE_OFN64405_a_in_3_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.634 36.957 35.662 37.12 ;
      END
   END FE_OFN64405_a_in_3_3

   PIN FE_OFN73421_n_32
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.33 0.0 49.358 0.163 ;
      END
   END FE_OFN73421_n_32

   PIN FE_OFN73591_n_44
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.274 36.957 36.302 37.12 ;
      END
   END FE_OFN73591_n_44

   PIN FE_OFN73647_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 2.29 57.728 2.318 ;
      END
   END FE_OFN73647_n_15

   PIN FE_OFN74017_n_31641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.565 2.162 57.728 2.19 ;
      END
   END FE_OFN74017_n_31641

   PIN FE_OFN74682_n_524
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 6.13 57.728 6.158 ;
      END
   END FE_OFN74682_n_524

   PIN FE_OFN85123_n_33
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.114 0.0 56.142 0.163 ;
      END
   END FE_OFN85123_n_33

   PIN FE_OFN85607_n_82
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.01 36.957 41.038 37.12 ;
      END
   END FE_OFN85607_n_82

   PIN FE_OFN85608_n_82
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.834 0.0 38.862 0.163 ;
      END
   END FE_OFN85608_n_82

   PIN FE_OFN86767_n_36757
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.898 0.163 22.926 ;
      END
   END FE_OFN86767_n_36757

   PIN FE_OFN91935_n_31635
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 2.354 57.728 2.382 ;
      END
   END FE_OFN91935_n_31635

   PIN FE_OFN91977_n_857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.106 36.957 45.134 37.12 ;
      END
   END FE_OFN91977_n_857

   PIN FE_OFN93495_ternarymux_ln49_0_unr61_z_9__4330986
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.482 0.163 26.51 ;
      END
   END FE_OFN93495_ternarymux_ln49_0_unr61_z_9__4330986

   PIN FE_OFN98121_n_32
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.138 36.957 57.166 37.12 ;
      END
   END FE_OFN98121_n_32

   PIN FE_RN_1501_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 5.938 57.728 5.966 ;
      END
   END FE_RN_1501_0

   PIN FE_RN_5563_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 19.122 57.728 19.15 ;
      END
   END FE_RN_5563_0

   PIN FE_RN_5983_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.93 0.163 18.958 ;
      END
   END FE_RN_5983_0

   PIN add_ln174_1_unr61_z_10__2985680
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.61 0.163 34.638 ;
      END
   END add_ln174_1_unr61_z_10__2985680

   PIN add_ln174_1_unr61_z_8__2227506
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.946 0.163 24.974 ;
      END
   END add_ln174_1_unr61_z_8__2227506

   PIN g2_m_82__5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 34.546 57.728 34.574 ;
      END
   END g2_m_82__5_

   PIN g2_q63_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 16.434 57.728 16.462 ;
      END
   END g2_q63_10_

   PIN g2_q63_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 34.61 57.728 34.638 ;
      END
   END g2_q63_11_

   PIN g2_q63_2__4327386
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 5.874 57.728 5.902 ;
      END
   END g2_q63_2__4327386

   PIN g2_q63_4__4327390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 2.482 57.728 2.51 ;
      END
   END g2_q63_4__4327390

   PIN g2_q63_6__4327379
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 22.898 57.728 22.926 ;
      END
   END g2_q63_6__4327379

   PIN g2_q63_7__4327380
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.098 36.957 50.126 37.12 ;
      END
   END g2_q63_7__4327380

   PIN g2_q63_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.218 36.957 47.246 37.12 ;
      END
   END g2_q63_9_

   PIN memread_edit_dist_g2_ln254_unr61_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 14.45 57.728 14.478 ;
      END
   END memread_edit_dist_g2_ln254_unr61_q_0_

   PIN memread_edit_dist_g2_ln254_unr61_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 4.658 57.728 4.686 ;
      END
   END memread_edit_dist_g2_ln254_unr61_q_1_

   PIN memread_edit_dist_g2_ln254_unr61_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 27.57 57.728 27.598 ;
      END
   END memread_edit_dist_g2_ln254_unr61_q_5_

   PIN memread_edit_dist_g2_ln254_unr61_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 18.802 57.728 18.83 ;
      END
   END memread_edit_dist_g2_ln254_unr61_q_8_

   PIN n_24340
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 10.674 57.728 10.702 ;
      END
   END n_24340

   PIN n_26697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.674 0.163 10.702 ;
      END
   END n_26697

   PIN n_27298
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 18.866 57.728 18.894 ;
      END
   END n_27298

   PIN n_27299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 25.074 57.728 25.102 ;
      END
   END n_27299

   PIN n_27447
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.802 0.082 10.83 ;
      END
   END n_27447

   PIN n_31764
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.346 0.0 55.374 0.163 ;
      END
   END n_31764

   PIN n_31953
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.914 36.957 36.942 37.12 ;
      END
   END n_31953

   PIN n_32018
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 16.306 57.728 16.334 ;
      END
   END n_32018

   PIN n_32973
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.762 36.957 35.79 37.12 ;
      END
   END n_32973

   PIN n_33099
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.162 36.957 50.19 37.12 ;
      END
   END n_33099

   PIN n_33228
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.682 0.163 21.71 ;
      END
   END n_33228

   PIN n_33242
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.514 0.163 30.542 ;
      END
   END n_33242

   PIN n_33306
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.546 0.163 34.574 ;
      END
   END n_33306

   PIN n_33604
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.178 0.163 16.206 ;
      END
   END n_33604

   PIN n_33628
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.026 0.163 31.054 ;
      END
   END n_33628

   PIN n_33629
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.482 0.163 34.51 ;
      END
   END n_33629

   PIN n_33671
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.994 0.163 19.022 ;
      END
   END n_33671

   PIN n_33727
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.962 0.163 22.99 ;
      END
   END n_33727

   PIN n_33944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.474 0.163 7.502 ;
      END
   END n_33944

   PIN n_34407
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.418 0.163 34.446 ;
      END
   END n_34407

   PIN n_35212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.626 0.082 24.654 ;
      END
   END n_35212

   PIN n_39172
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.546 0.163 10.574 ;
      END
   END n_39172

   PIN n_39327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.61 0.163 10.638 ;
      END
   END n_39327

   PIN n_39343
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.578 0.163 14.606 ;
      END
   END n_39343

   PIN n_39370
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.106 0.163 13.134 ;
      END
   END n_39370

   PIN n_43334
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.946 0.0 24.974 0.163 ;
      END
   END n_43334

   PIN n_60455
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.818 0.0 32.846 0.163 ;
      END
   END n_60455

   PIN n_60469
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 1.714 57.728 1.742 ;
      END
   END n_60469

   PIN n_60475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 24.69 57.728 24.718 ;
      END
   END n_60475

   PIN n_60667
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 1.778 57.728 1.806 ;
      END
   END n_60667

   PIN n_64828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.646 24.818 57.728 24.846 ;
      END
   END n_64828

   PIN n_66478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.306 0.163 16.334 ;
      END
   END n_66478

   PIN ternarymux_ln49_0_unr61_z_8__4330990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.338 0.0 36.366 0.163 ;
      END
   END ternarymux_ln49_0_unr61_z_8__4330990

   PIN ternarymux_ln49_0_unr62_z_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.594 0.163 4.622 ;
      END
   END ternarymux_ln49_0_unr62_z_1_

   PIN ternarymux_ln49_0_unr62_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.922 0.163 15.95 ;
      END
   END ternarymux_ln49_0_unr62_z_3_

   PIN ternarymux_ln49_0_unr62_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.05 0.163 16.078 ;
      END
   END ternarymux_ln49_0_unr62_z_4_

   PIN ternarymux_ln49_0_unr62_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.802 0.163 18.83 ;
      END
   END ternarymux_ln49_0_unr62_z_5_

   PIN ternarymux_ln49_0_unr62_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.114 0.163 16.142 ;
      END
   END ternarymux_ln49_0_unr62_z_7_

   PIN ternarymux_ln49_0_unr82_z_10__4331318
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.354 0.163 34.382 ;
      END
   END ternarymux_ln49_0_unr82_z_10__4331318

   PIN ternarymux_ln49_0_unr82_z_8__4331326
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 16.37 57.728 16.398 ;
      END
   END ternarymux_ln49_0_unr82_z_8__4331326

   PIN ternarymux_ln49_5_unr62_z_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.754 0.163 24.782 ;
      END
   END ternarymux_ln49_5_unr62_z_0_

   PIN ternarymux_ln49_6_unr82_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 14.514 57.728 14.542 ;
      END
   END ternarymux_ln49_6_unr82_z_12_

   PIN ternarymux_ln49_8_unr82_z_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 21.682 57.728 21.71 ;
      END
   END ternarymux_ln49_8_unr82_z_11_

   PIN FE_OCPN57527_FE_OFN47118_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 10.61 57.728 10.638 ;
      END
   END FE_OCPN57527_FE_OFN47118_n_23039

   PIN FE_OCPN57867_n_93
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 14.386 57.728 14.414 ;
      END
   END FE_OCPN57867_n_93

   PIN FE_OCPN58733_FE_OFN46361_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.498 36.957 48.526 37.12 ;
      END
   END FE_OCPN58733_FE_OFN46361_n_67216

   PIN FE_OCPN60536_FE_OFN48705_n_59125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.442 0.0 43.47 0.163 ;
      END
   END FE_OCPN60536_FE_OFN48705_n_59125

   PIN FE_OCPN62476_n_65256
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.058 36.957 19.086 37.12 ;
      END
   END FE_OCPN62476_n_65256

   PIN FE_OCPN78686_ternarymux_ln49_0_unr62_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.77 0.163 22.798 ;
      END
   END FE_OCPN78686_ternarymux_ln49_0_unr62_z_4_

   PIN FE_OCPN78960_add_ln174_1_unr81_z_8__2227792
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 26.802 57.728 26.83 ;
      END
   END FE_OCPN78960_add_ln174_1_unr81_z_8__2227792

   PIN FE_OCP_DRV_N76505_n_32047
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 18.93 57.728 18.958 ;
      END
   END FE_OCP_DRV_N76505_n_32047

   PIN FE_OFN29317_n_524
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.082 0.0 4.11 0.163 ;
      END
   END FE_OFN29317_n_524

   PIN FE_OFN30108_n_36239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 15.922 57.728 15.95 ;
      END
   END FE_OFN30108_n_36239

   PIN FE_OFN30153_n_36584
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 14.322 57.728 14.35 ;
      END
   END FE_OFN30153_n_36584

   PIN FE_OFN30155_n_36438
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.282 0.0 47.31 0.163 ;
      END
   END FE_OFN30155_n_36438

   PIN FE_OFN30163_n_36334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 6.642 57.728 6.67 ;
      END
   END FE_OFN30163_n_36334

   PIN FE_OFN30326_n_36003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 7.41 57.728 7.438 ;
      END
   END FE_OFN30326_n_36003

   PIN FE_OFN30400_n_35970
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 10.546 57.728 10.574 ;
      END
   END FE_OFN30400_n_35970

   PIN FE_OFN30637_n_36637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 16.242 57.728 16.27 ;
      END
   END FE_OFN30637_n_36637

   PIN FE_OFN30801_n_36371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 2.162 57.728 2.19 ;
      END
   END FE_OFN30801_n_36371

   PIN FE_OFN31996_n_31637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 27.122 0.163 27.15 ;
      END
   END FE_OFN31996_n_31637

   PIN FE_OFN34194_n_82
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.042 36.957 53.07 37.12 ;
      END
   END FE_OFN34194_n_82

   PIN FE_OFN42374_n_44
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.338 0.0 36.366 0.163 ;
      END
   END FE_OFN42374_n_44

   PIN FE_OFN42487_n_33
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.73 36.957 47.758 37.12 ;
      END
   END FE_OFN42487_n_33

   PIN FE_OFN46247_a_in_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.514 0.163 14.542 ;
      END
   END FE_OFN46247_a_in_6_2

   PIN FE_OFN46272_a_in_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.698 36.957 35.726 37.12 ;
      END
   END FE_OFN46272_a_in_3_3

   PIN FE_OFN47675_n_22885
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.794 0.0 55.822 0.163 ;
      END
   END FE_OFN47675_n_22885

   PIN FE_OFN47898_n_31635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.162 0.163 2.19 ;
      END
   END FE_OFN47898_n_31635

   PIN FE_OFN48370_n_31641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.578 0.163 30.606 ;
      END
   END FE_OFN48370_n_31641

   PIN FE_OFN50337_n_64841
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.962 0.163 30.99 ;
      END
   END FE_OFN50337_n_64841

   PIN FE_OFN50338_n_64841
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 16.114 0.163 16.142 ;
      END
   END FE_OFN50338_n_64841

   PIN FE_OFN50556_lt_ln49_6_unr82_z
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.646 10.802 57.728 10.83 ;
      END
   END FE_OFN50556_lt_ln49_6_unr82_z

   PIN FE_OFN50580_lt_ln49_6_unr61_z
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.642 0.082 22.67 ;
      END
   END FE_OFN50580_lt_ln49_6_unr61_z

   PIN FE_OFN53691_n_91
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.962 0.0 6.99 0.163 ;
      END
   END FE_OFN53691_n_91

   PIN FE_OFN55966_ternarymux_ln49_0_unr61_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 57.565 1.714 57.728 1.742 ;
      END
   END FE_OFN55966_ternarymux_ln49_0_unr61_z_5_

   PIN FE_OFN55978_ternarymux_ln49_0_unr61_z_10__4330982
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.746 0.0 53.774 0.163 ;
      END
   END FE_OFN55978_ternarymux_ln49_0_unr61_z_10__4330982

   PIN FE_OFN70914_memwrite_edit_dist_g2_ln280_unr61_en_0__4469706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.194 36.957 14.222 37.12 ;
      END
   END FE_OFN70914_memwrite_edit_dist_g2_ln280_unr61_en_0__4469706

   PIN FE_OFN70915_n_21264
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.714 36.957 17.742 37.12 ;
      END
   END FE_OFN70915_n_21264

   PIN FE_OFN85983_FE_OCPN60599_FE_OFN48344_n_31639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.346 0.163 31.374 ;
      END
   END FE_OFN85983_FE_OCPN60599_FE_OFN48344_n_31639

   PIN FE_OFN86656_n_36241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 13.106 57.728 13.134 ;
      END
   END FE_OFN86656_n_36241

   PIN FE_OFN86766_n_36757
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 16.178 57.728 16.206 ;
      END
   END FE_OFN86766_n_36757

   PIN FE_OFN88247_n_31634
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 4.722 57.728 4.75 ;
      END
   END FE_OFN88247_n_31634

   PIN FE_OFN90783_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 10.482 57.728 10.51 ;
      END
   END FE_OFN90783_n_67217

   PIN FE_OFN91976_n_857
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.618 0.0 45.646 0.163 ;
      END
   END FE_OFN91976_n_857

   PIN FE_OFN92515_n_31642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.474 36.957 15.502 37.12 ;
      END
   END FE_OFN92515_n_31642

   PIN FE_OFN93183_FE_OCPN61464_FE_OFN48299_n_31625
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.522 36.957 41.55 37.12 ;
      END
   END FE_OFN93183_FE_OCPN61464_FE_OFN48299_n_31625

   PIN FE_OFN98340_ternarymux_ln49_0_unr62_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.482 0.163 18.51 ;
      END
   END FE_OFN98340_ternarymux_ln49_0_unr62_z_2_

   PIN FE_RN_1499_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.914 0.0 52.942 0.163 ;
      END
   END FE_RN_1499_0

   PIN a_in_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.634 0.163 27.662 ;
      END
   END a_in_3_3

   PIN add_ln174_1_unr60_z_10__2985662
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.05 0.0 56.078 0.163 ;
      END
   END add_ln174_1_unr60_z_10__2985662

   PIN add_ln174_1_unr60_z_8__2227484
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.922 0.0 55.95 0.163 ;
      END
   END add_ln174_1_unr60_z_8__2227484

   PIN add_ln174_1_unr60_z_9__2985661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.986 0.0 56.014 0.163 ;
      END
   END add_ln174_1_unr60_z_9__2985661

   PIN add_ln174_1_unr81_z_10__2985914
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.33 36.957 49.358 37.12 ;
      END
   END add_ln174_1_unr81_z_10__2985914

   PIN add_ln174_1_unr81_z_9__2985913
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 31.09 57.728 31.118 ;
      END
   END add_ln174_1_unr81_z_9__2985913

   PIN g2_m_81__6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.642 0.163 30.67 ;
      END
   END g2_m_81__6_

   PIN g2_q63_3__4327387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.858 0.0 47.886 0.163 ;
      END
   END g2_q63_3__4327387

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.906 0.0 41.934 0.082 ;
      END
   END ispd_clk

   PIN memread_edit_dist_a_ln268_unr124_a_33__4330321
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.082 0.0 4.11 0.163 ;
      END
   END memread_edit_dist_a_ln268_unr124_a_33__4330321

   PIN mux_g_ln477_q_538_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.106 36.957 53.134 37.12 ;
      END
   END mux_g_ln477_q_538_

   PIN n_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.482 0.0 18.51 0.163 ;
      END
   END n_15

   PIN n_26724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 24.626 57.728 24.654 ;
      END
   END n_26724

   PIN n_27093
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.482 0.163 10.51 ;
      END
   END n_27093

   PIN n_27289
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 24.562 57.728 24.59 ;
      END
   END n_27289

   PIN n_27691
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.098 0.0 34.126 0.163 ;
      END
   END n_27691

   PIN n_28399
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.646 30.962 57.728 30.99 ;
      END
   END n_28399

   PIN n_28421
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 21.81 57.728 21.838 ;
      END
   END n_28421

   PIN n_28422
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 22.834 57.728 22.862 ;
      END
   END n_28422

   PIN n_28515
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 22.77 57.728 22.798 ;
      END
   END n_28515

   PIN n_2966
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.858 36.957 47.886 37.12 ;
      END
   END n_2966

   PIN n_31796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.042 36.957 45.07 37.12 ;
      END
   END n_31796

   PIN n_32
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.402 0.0 44.43 0.163 ;
      END
   END n_32

   PIN n_33098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.162 36.957 50.19 37.12 ;
      END
   END n_33098

   PIN n_33248
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.354 0.0 26.382 0.163 ;
      END
   END n_33248

   PIN n_33317
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 19.058 57.728 19.086 ;
      END
   END n_33317

   PIN n_33768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.018 0.0 36.046 0.163 ;
      END
   END n_33768

   PIN n_34371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 15.986 0.163 16.014 ;
      END
   END n_34371

   PIN n_35200
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.466 0.0 20.494 0.163 ;
      END
   END n_35200

   PIN n_35944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 18.994 57.728 19.022 ;
      END
   END n_35944

   PIN n_36245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 4.594 57.728 4.622 ;
      END
   END n_36245

   PIN n_39238
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.754 0.163 24.782 ;
      END
   END n_39238

   PIN n_48546
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.646 16.05 57.728 16.078 ;
      END
   END n_48546

   PIN n_51746
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.45 0.163 14.478 ;
      END
   END n_51746

   PIN n_59964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.646 22.642 57.728 22.67 ;
      END
   END n_59964

   PIN n_60462
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.874 0.163 5.902 ;
      END
   END n_60462

   PIN n_60666
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 27.122 57.728 27.15 ;
      END
   END n_60666

   PIN n_61220
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 25.01 57.728 25.038 ;
      END
   END n_61220

   PIN n_61225
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 21.618 57.728 21.646 ;
      END
   END n_61225

   PIN n_62440
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.386 0.163 14.414 ;
      END
   END n_62440

   PIN n_62441
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.322 0.163 14.35 ;
      END
   END n_62441

   PIN n_62442
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.938 0.163 5.966 ;
      END
   END n_62442

   PIN n_62443
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.242 0.0 24.27 0.163 ;
      END
   END n_62443

   PIN n_64842
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 22.962 57.728 22.99 ;
      END
   END n_64842

   PIN n_66477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.234 0.0 53.262 0.163 ;
      END
   END n_66477

   PIN ternarymux_ln49_0_unr61_z_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.65 0.0 33.678 0.163 ;
      END
   END ternarymux_ln49_0_unr61_z_0_

   PIN ternarymux_ln49_0_unr61_z_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.738 0.0 18.766 0.163 ;
      END
   END ternarymux_ln49_0_unr61_z_1_

   PIN ternarymux_ln49_0_unr61_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.194 0.0 30.222 0.163 ;
      END
   END ternarymux_ln49_0_unr61_z_2_

   PIN ternarymux_ln49_0_unr61_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.394 0.0 17.422 0.163 ;
      END
   END ternarymux_ln49_0_unr61_z_3_

   PIN ternarymux_ln49_0_unr61_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END ternarymux_ln49_0_unr61_z_4_

   PIN ternarymux_ln49_0_unr61_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.578 0.0 22.606 0.163 ;
      END
   END ternarymux_ln49_0_unr61_z_6_

   PIN ternarymux_ln49_0_unr61_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.002 0.0 14.03 0.163 ;
      END
   END ternarymux_ln49_0_unr61_z_7_

   PIN ternarymux_ln49_0_unr61_z_9__4330986
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.754 0.0 40.782 0.163 ;
      END
   END ternarymux_ln49_0_unr61_z_9__4330986

   PIN ternarymux_ln49_0_unr62_z_8__4331006
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.802 0.163 18.83 ;
      END
   END ternarymux_ln49_0_unr62_z_8__4331006

   PIN ternarymux_ln49_0_unr62_z_9__4331002
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.546 0.163 26.574 ;
      END
   END ternarymux_ln49_0_unr62_z_9__4331002

   PIN ternarymux_ln49_0_unr82_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 24.946 57.728 24.974 ;
      END
   END ternarymux_ln49_0_unr82_z_3_

   PIN ternarymux_ln49_0_unr82_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 34.482 57.728 34.51 ;
      END
   END ternarymux_ln49_0_unr82_z_5_

   PIN ternarymux_ln49_8_unr82_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 57.565 21.746 57.728 21.774 ;
      END
   END ternarymux_ln49_8_unr82_z_9_

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 57.728 37.12 ;
      LAYER V1 ;
         RECT 0.0 0.0 57.728 37.12 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 57.728 37.12 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 57.728 37.12 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 57.728 37.12 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 57.728 37.12 ;
      LAYER M1 ;
         RECT 0.0 0.0 57.728 37.12 ;
   END
END h2_mgc_edit_dist_a

MACRO h1_mgc_edit_dist_a
   CLASS BLOCK ;
   FOREIGN h1 ;
   ORIGIN 0 0 ;
   SIZE 58.56 BY 80.0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN56133_n_35331
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 54.322 58.56 54.35 ;
      END
   END FE_OCPN56133_n_35331

   PIN FE_OCPN57867_n_93
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.946 0.0 56.974 0.163 ;
      END
   END FE_OCPN57867_n_93

   PIN FE_OCPN58711_n_33467_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.442 0.0 35.47 0.163 ;
      END
   END FE_OCPN58711_n_33467_bar

   PIN FE_OCPN60456_memread_edit_dist_a_ln268_unr124_a_9__4329837
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 17.522 58.56 17.55 ;
      END
   END FE_OCPN60456_memread_edit_dist_a_ln268_unr124_a_9__4329837

   PIN FE_OCPN60530_FE_OFN48705_n_59125
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.458 0.0 9.486 0.163 ;
      END
   END FE_OCPN60530_FE_OFN48705_n_59125

   PIN FE_OCPN61465_FE_OFN48299_n_31625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 46.066 0.163 46.094 ;
      END
   END FE_OCPN61465_FE_OFN48299_n_31625

   PIN FE_OCPN62334_n_58046
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.834 0.163 62.862 ;
      END
   END FE_OCPN62334_n_58046

   PIN FE_OCPN62350_n_65199
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.506 0.0 43.534 0.163 ;
      END
   END FE_OCPN62350_n_65199

   PIN FE_OCPN62854_n_33487_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.754 0.0 40.782 0.163 ;
      END
   END FE_OCPN62854_n_33487_bar

   PIN FE_OCPN63056_FE_OFN47982_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 20.018 58.56 20.046 ;
      END
   END FE_OCPN63056_FE_OFN47982_n_23035

   PIN FE_OCPN63788_FE_OFN48830_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.162 0.0 18.19 0.163 ;
      END
   END FE_OCPN63788_FE_OFN48830_n_31626

   PIN FE_OCPN63795_FE_OFN48307_n_31634
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.402 0.0 12.43 0.163 ;
      END
   END FE_OCPN63795_FE_OFN48307_n_31634

   PIN FE_OCPN78052_FE_OFN48367_n_31641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.25 0.163 75.278 ;
      END
   END FE_OCPN78052_FE_OFN48367_n_31641

   PIN FE_OCPN95861_n_58050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.162 79.837 18.19 80.0 ;
      END
   END FE_OCPN95861_n_58050

   PIN FE_OFN28637_n_36328
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 45.81 58.56 45.838 ;
      END
   END FE_OFN28637_n_36328

   PIN FE_OFN28734_n_40187
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.642 0.0 6.67 0.082 ;
      END
   END FE_OFN28734_n_40187

   PIN FE_OFN30022_n_36839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 66.098 0.163 66.126 ;
      END
   END FE_OFN30022_n_36839

   PIN FE_OFN30049_n_36035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.442 0.163 35.47 ;
      END
   END FE_OFN30049_n_36035

   PIN FE_OFN30051_n_36014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.714 0.163 57.742 ;
      END
   END FE_OFN30051_n_36014

   PIN FE_OFN30065_n_37068
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.986 0.163 64.014 ;
      END
   END FE_OFN30065_n_37068

   PIN FE_OFN30075_n_36916
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 42.93 0.163 42.958 ;
      END
   END FE_OFN30075_n_36916

   PIN FE_OFN30206_n_36803
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.842 0.163 25.87 ;
      END
   END FE_OFN30206_n_36803

   PIN FE_OFN30245_n_37046
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 51.57 0.163 51.598 ;
      END
   END FE_OFN30245_n_37046

   PIN FE_OFN30248_n_37029
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.282 0.163 31.31 ;
      END
   END FE_OFN30248_n_37029

   PIN FE_OFN30266_n_36785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.802 0.163 42.83 ;
      END
   END FE_OFN30266_n_36785

   PIN FE_OFN30301_n_36379
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 17.01 0.163 17.038 ;
      END
   END FE_OFN30301_n_36379

   PIN FE_OFN30337_n_36733
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 51.634 0.163 51.662 ;
      END
   END FE_OFN30337_n_36733

   PIN FE_OFN30356_n_35984
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 65.97 0.163 65.998 ;
      END
   END FE_OFN30356_n_35984

   PIN FE_OFN30389_n_34771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.754 0.0 56.782 0.163 ;
      END
   END FE_OFN30389_n_34771

   PIN FE_OFN30460_n_36563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.562 0.163 48.59 ;
      END
   END FE_OFN30460_n_36563

   PIN FE_OFN30471_n_35975
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 70.642 0.163 70.67 ;
      END
   END FE_OFN30471_n_35975

   PIN FE_OFN30521_n_36965
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.482 0.163 26.51 ;
      END
   END FE_OFN30521_n_36965

   PIN FE_OFN30531_n_36390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.33 0.163 57.358 ;
      END
   END FE_OFN30531_n_36390

   PIN FE_OFN30574_n_36953
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.082 0.163 60.11 ;
      END
   END FE_OFN30574_n_36953

   PIN FE_OFN30590_n_36899
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.986 0.163 40.014 ;
      END
   END FE_OFN30590_n_36899

   PIN FE_OFN30594_n_36874
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.354 0.163 34.382 ;
      END
   END FE_OFN30594_n_36874

   PIN FE_OFN30641_n_36622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 42.994 0.163 43.022 ;
      END
   END FE_OFN30641_n_36622

   PIN FE_OFN30660_n_36401
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.85 0.163 68.878 ;
      END
   END FE_OFN30660_n_36401

   PIN FE_OFN30662_n_36399
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 66.034 0.163 66.062 ;
      END
   END FE_OFN30662_n_36399

   PIN FE_OFN30685_n_36201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 29.042 0.163 29.07 ;
      END
   END FE_OFN30685_n_36201

   PIN FE_OFN30698_n_36086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.994 0.163 35.022 ;
      END
   END FE_OFN30698_n_36086

   PIN FE_OFN30707_n_36073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.866 0.163 42.894 ;
      END
   END FE_OFN30707_n_36073

   PIN FE_OFN30717_n_36030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.666 0.163 31.694 ;
      END
   END FE_OFN30717_n_36030

   PIN FE_OFN30724_n_36015
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 55.026 0.163 55.054 ;
      END
   END FE_OFN30724_n_36015

   PIN FE_OFN30729_n_35986
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.282 0.163 23.31 ;
      END
   END FE_OFN30729_n_35986

   PIN FE_OFN30733_n_35978
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.562 0.163 72.59 ;
      END
   END FE_OFN30733_n_35978

   PIN FE_OFN30796_n_36565
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.01 0.163 33.038 ;
      END
   END FE_OFN30796_n_36565

   PIN FE_OFN30810_n_34732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.57 0.0 35.598 0.163 ;
      END
   END FE_OFN30810_n_34732

   PIN FE_OFN30812_n_34732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 34.29 58.56 34.318 ;
      END
   END FE_OFN30812_n_34732

   PIN FE_OFN30828_n_36787
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.098 79.837 26.126 80.0 ;
      END
   END FE_OFN30828_n_36787

   PIN FE_OFN30862_n_34779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.626 0.0 32.654 0.163 ;
      END
   END FE_OFN30862_n_34779

   PIN FE_OFN30869_n_36922
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 78.322 0.163 78.35 ;
      END
   END FE_OFN30869_n_36922

   PIN FE_OFN30904_n_35995
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.93 0.163 42.958 ;
      END
   END FE_OFN30904_n_35995

   PIN FE_OFN31034_n_34785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.186 0.0 51.214 0.163 ;
      END
   END FE_OFN31034_n_34785

   PIN FE_OFN32007_n_31638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.058 0.163 43.086 ;
      END
   END FE_OFN32007_n_31638

   PIN FE_OFN32021_n_31639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.002 0.163 14.03 ;
      END
   END FE_OFN32021_n_31639

   PIN FE_OFN32360_n_21259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.57 0.163 51.598 ;
      END
   END FE_OFN32360_n_21259

   PIN FE_OFN33793_n_3370
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.562 0.0 32.59 0.163 ;
      END
   END FE_OFN33793_n_3370

   PIN FE_OFN34105_n_86
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.69 0.0 16.718 0.163 ;
      END
   END FE_OFN34105_n_86

   PIN FE_OFN34914_n_53413
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.626 0.163 48.654 ;
      END
   END FE_OFN34914_n_53413

   PIN FE_OFN34942_n_51091
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.698 0.163 51.726 ;
      END
   END FE_OFN34942_n_51091

   PIN FE_OFN41931_n_230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.082 0.0 44.11 0.163 ;
      END
   END FE_OFN41931_n_230

   PIN FE_OFN42169_n_53
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.602 79.837 55.63 80.0 ;
      END
   END FE_OFN42169_n_53

   PIN FE_OFN42913_n_3242
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 55.858 58.56 55.886 ;
      END
   END FE_OFN42913_n_3242

   PIN FE_OFN43005_n_35325
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.538 0.0 55.566 0.163 ;
      END
   END FE_OFN43005_n_35325

   PIN FE_OFN43958_mux_g_ln477_q_520_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.986 79.837 40.014 80.0 ;
      END
   END FE_OFN43958_mux_g_ln477_q_520_

   PIN FE_OFN47854_n_23045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.65 79.837 33.678 80.0 ;
      END
   END FE_OFN47854_n_23045

   PIN FE_OFN48299_n_31625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.866 0.0 26.894 0.163 ;
      END
   END FE_OFN48299_n_31625

   PIN FE_OFN48313_n_31634
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.202 0.082 57.23 ;
      END
   END FE_OFN48313_n_31634

   PIN FE_OFN48316_n_31634
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.322 0.163 46.35 ;
      END
   END FE_OFN48316_n_31634

   PIN FE_OFN48344_n_31639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.762 0.0 3.79 0.163 ;
      END
   END FE_OFN48344_n_31639

   PIN FE_OFN48367_n_31641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.298 0.163 37.326 ;
      END
   END FE_OFN48367_n_31641

   PIN FE_OFN48368_n_31641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.418 0.0 2.446 0.163 ;
      END
   END FE_OFN48368_n_31641

   PIN FE_OFN48708_n_59125
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.042 0.163 37.07 ;
      END
   END FE_OFN48708_n_59125

   PIN FE_OFN48845_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.106 0.163 37.134 ;
      END
   END FE_OFN48845_n_31626

   PIN FE_OFN48846_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.674 0.163 74.702 ;
      END
   END FE_OFN48846_n_31626

   PIN FE_OFN48848_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.834 0.0 46.862 0.163 ;
      END
   END FE_OFN48848_n_31626

   PIN FE_OFN49702_n_87
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.226 79.837 18.254 80.0 ;
      END
   END FE_OFN49702_n_87

   PIN FE_OFN49703_n_87
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.746 79.837 29.774 80.0 ;
      END
   END FE_OFN49703_n_87

   PIN FE_OFN50544_lt_ln49_6_unr75_z
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.586 0.163 57.614 ;
      END
   END FE_OFN50544_lt_ln49_6_unr75_z

   PIN FE_OFN50546_lt_ln49_6_unr75_z
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.002 0.163 54.03 ;
      END
   END FE_OFN50546_lt_ln49_6_unr75_z

   PIN FE_OFN70357_n_36808
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 69.426 58.56 69.454 ;
      END
   END FE_OFN70357_n_36808

   PIN FE_OFN71105_memwrite_edit_dist_g2_ln280_unr73_en_0__4469519
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 74.674 0.163 74.702 ;
      END
   END FE_OFN71105_memwrite_edit_dist_g2_ln280_unr73_en_0__4469519

   PIN FE_OFN71827_n_51730
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.714 0.163 65.742 ;
      END
   END FE_OFN71827_n_51730

   PIN FE_OFN73372_n_20
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.378 79.837 51.406 80.0 ;
      END
   END FE_OFN73372_n_20

   PIN FE_OFN73646_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.802 79.837 34.83 80.0 ;
      END
   END FE_OFN73646_n_15

   PIN FE_OFN73661_n_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.042 79.837 21.07 80.0 ;
      END
   END FE_OFN73661_n_29

   PIN FE_OFN73975_n_32261
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.362 0.163 53.39 ;
      END
   END FE_OFN73975_n_32261

   PIN FE_OFN74037_n_31638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.802 0.0 26.83 0.163 ;
      END
   END FE_OFN74037_n_31638

   PIN FE_OFN74082_n_59052
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.818 0.163 16.846 ;
      END
   END FE_OFN74082_n_59052

   PIN FE_OFN74310_n_61
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 1.586 58.56 1.614 ;
      END
   END FE_OFN74310_n_61

   PIN FE_OFN74580_n_79
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.226 0.0 18.254 0.163 ;
      END
   END FE_OFN74580_n_79

   PIN FE_OFN74879_n_36980
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 19.954 0.163 19.982 ;
      END
   END FE_OFN74879_n_36980

   PIN FE_OFN74969_n_36218
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.922 0.163 23.95 ;
      END
   END FE_OFN74969_n_36218

   PIN FE_OFN75080_n_34770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.946 0.0 56.974 0.163 ;
      END
   END FE_OFN75080_n_34770

   PIN FE_OFN75216_n_35297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.898 79.837 46.926 80.0 ;
      END
   END FE_OFN75216_n_35297

   PIN FE_OFN75258_n_35301
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 4.85 58.56 4.878 ;
      END
   END FE_OFN75258_n_35301

   PIN FE_OFN75313_n_35325
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 45.938 58.56 45.966 ;
      END
   END FE_OFN75313_n_35325

   PIN FE_OFN75550_FE_OCPN62021_FE_OFN50813_n_67216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 5.81 58.56 5.838 ;
      END
   END FE_OFN75550_FE_OCPN62021_FE_OFN50813_n_67216

   PIN FE_OFN75725_n_35331
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 78.386 58.56 78.414 ;
      END
   END FE_OFN75725_n_35331

   PIN FE_OFN84025_n_21287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.17 0.163 37.198 ;
      END
   END FE_OFN84025_n_21287

   PIN FE_OFN84037_n_7936
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 8.626 58.56 8.654 ;
      END
   END FE_OFN84037_n_7936

   PIN FE_OFN85021_n_57
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.602 79.837 47.63 80.0 ;
      END
   END FE_OFN85021_n_57

   PIN FE_OFN85096_n_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.922 79.837 23.95 80.0 ;
      END
   END FE_OFN85096_n_30

   PIN FE_OFN85107_n_53
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.682 79.837 45.71 80.0 ;
      END
   END FE_OFN85107_n_53

   PIN FE_OFN85118_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 75.762 58.56 75.79 ;
      END
   END FE_OFN85118_n_15

   PIN FE_OFN85990_n_31637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.106 0.163 45.134 ;
      END
   END FE_OFN85990_n_31637

   PIN FE_OFN86082_g2_q72_2__4327665
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 28.53 58.56 28.558 ;
      END
   END FE_OFN86082_g2_q72_2__4327665

   PIN FE_OFN86624_n_36643
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.586 0.163 49.614 ;
      END
   END FE_OFN86624_n_36643

   PIN FE_OFN86680_n_36864
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.818 0.163 48.846 ;
      END
   END FE_OFN86680_n_36864

   PIN FE_OFN86686_n_35998
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 23.666 0.163 23.694 ;
      END
   END FE_OFN86686_n_35998

   PIN FE_OFN86751_n_36820
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.634 0.163 51.662 ;
      END
   END FE_OFN86751_n_36820

   PIN FE_OFN86757_n_36061
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.346 0.163 31.374 ;
      END
   END FE_OFN86757_n_36061

   PIN FE_OFN86879_n_36948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 15.73 0.163 15.758 ;
      END
   END FE_OFN86879_n_36948

   PIN FE_OFN86936_n_36221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.554 0.163 77.582 ;
      END
   END FE_OFN86936_n_36221

   PIN FE_OFN87036_n_35936
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.418 0.163 34.446 ;
      END
   END FE_OFN87036_n_35936

   PIN FE_OFN87056_n_36888
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.778 0.163 57.806 ;
      END
   END FE_OFN87056_n_36888

   PIN FE_OFN87975_n_35283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 23.282 58.56 23.31 ;
      END
   END FE_OFN87975_n_35283

   PIN FE_OFN88306_n_65239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.642 0.163 54.67 ;
      END
   END FE_OFN88306_n_65239

   PIN FE_OFN94568_n_31625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.826 0.0 19.854 0.163 ;
      END
   END FE_OFN94568_n_31625

   PIN FE_OFN94908_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 1.522 58.56 1.55 ;
      END
   END FE_OFN94908_n_31626

   PIN FE_OFN95909_n_65250
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.05 0.163 40.078 ;
      END
   END FE_OFN95909_n_65250

   PIN FE_OFN98159_n_230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.594 79.837 52.622 80.0 ;
      END
   END FE_OFN98159_n_230

   PIN FE_OFN98509_n_37004
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 51.698 0.163 51.726 ;
      END
   END FE_OFN98509_n_37004

   PIN FE_OFN98531_n_36062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.25 0.163 27.278 ;
      END
   END FE_OFN98531_n_36062

   PIN FE_RN_3498_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.85 0.163 68.878 ;
      END
   END FE_RN_3498_0

   PIN add_85532_72_n_4327722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 69.362 0.163 69.39 ;
      END
   END add_85532_72_n_4327722

   PIN add_85538_72_n_4327812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.554 0.0 29.582 0.163 ;
      END
   END add_85538_72_n_4327812

   PIN g2_bridge202_rtl_ce_en_3755253_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.17 0.082 69.198 ;
      END
   END g2_bridge202_rtl_ce_en_3755253_bar

   PIN g2_bridge208_rtl_ce_en_3756288
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.81 0.163 13.838 ;
      END
   END g2_bridge208_rtl_ce_en_3756288

   PIN g2_q72_1__4327663
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.866 0.163 34.894 ;
      END
   END g2_q72_1__4327663

   PIN g2_q77_1__4327814
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 19.89 58.56 19.918 ;
      END
   END g2_q77_1__4327814

   PIN g2_q77_3__4327817
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 23.026 58.56 23.054 ;
      END
   END g2_q77_3__4327817

   PIN g2_q78_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.114 0.0 32.142 0.163 ;
      END
   END g2_q78_10_

   PIN g2_q78_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.322 0.0 38.35 0.163 ;
      END
   END g2_q78_8_

   PIN gt_93966_62_n_89
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.202 0.163 17.23 ;
      END
   END gt_93966_62_n_89

   PIN memread_edit_dist_a_ln268_unr124_a_21__4330189
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 30.386 58.56 30.414 ;
      END
   END memread_edit_dist_a_ln268_unr124_a_21__4330189

   PIN memread_edit_dist_g2_ln254_unr67_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 8.37 58.56 8.398 ;
      END
   END memread_edit_dist_g2_ln254_unr67_q_10_

   PIN memread_edit_dist_g2_ln254_unr67_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.498 0.0 56.526 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr67_q_1_

   PIN memread_edit_dist_g2_ln254_unr67_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.962 58.56 22.99 ;
      END
   END memread_edit_dist_g2_ln254_unr67_q_5_

   PIN memread_edit_dist_g2_ln254_unr68_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.618 0.0 29.646 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_10_

   PIN memread_edit_dist_g2_ln254_unr68_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.178 0.0 56.206 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_3_

   PIN memread_edit_dist_g2_ln254_unr69_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 11.378 58.56 11.406 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_4_

   PIN memread_edit_dist_g2_ln254_unr70_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 35.506 58.56 35.534 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_0_

   PIN memread_edit_dist_g2_ln254_unr70_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.498 0.0 40.526 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_10_

   PIN memread_edit_dist_g2_ln254_unr70_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 4.914 58.56 4.942 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_1_

   PIN memread_edit_dist_g2_ln254_unr70_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 2.738 58.56 2.766 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_3_

   PIN memread_edit_dist_g2_ln254_unr70_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 11.442 58.56 11.47 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_5_

   PIN memread_edit_dist_g2_ln254_unr70_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 29.746 58.56 29.774 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_7_

   PIN memread_edit_dist_g2_ln254_unr71_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 42.93 58.56 42.958 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_0_

   PIN memread_edit_dist_g2_ln254_unr71_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 2.802 58.56 2.83 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_1_

   PIN memread_edit_dist_g2_ln254_unr71_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 25.714 58.56 25.742 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_2_

   PIN memread_edit_dist_g2_ln254_unr71_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 54.514 58.56 54.542 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_3_

   PIN memread_edit_dist_g2_ln254_unr71_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 40.562 58.56 40.59 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_5_

   PIN memread_edit_dist_g2_ln254_unr71_q_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 14.066 58.56 14.094 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_6_

   PIN memread_edit_dist_g2_ln254_unr71_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 17.074 58.56 17.102 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_7_

   PIN memread_edit_dist_g2_ln254_unr72_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 39.986 58.56 40.014 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_0_

   PIN memread_edit_dist_g2_ln254_unr72_q_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 17.138 58.56 17.166 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_11_

   PIN memread_edit_dist_g2_ln254_unr72_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.786 0.0 52.814 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_1_

   PIN memread_edit_dist_g2_ln254_unr72_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 17.202 58.56 17.23 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_2_

   PIN memread_edit_dist_g2_ln254_unr72_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 54.578 58.56 54.606 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_3_

   PIN memread_edit_dist_g2_ln254_unr72_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 46.002 58.56 46.03 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_4_

   PIN memread_edit_dist_g2_ln254_unr72_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 57.394 58.56 57.422 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_5_

   PIN memread_edit_dist_g2_ln254_unr76_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.05 0.0 40.078 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_0_

   PIN memread_edit_dist_g2_ln254_unr76_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.698 0.0 43.726 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_1_

   PIN memread_edit_dist_g2_ln254_unr76_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.298 0.0 45.326 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_2_

   PIN memread_edit_dist_g2_ln254_unr76_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 49.714 0.0 49.742 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_3_

   PIN memread_edit_dist_g2_ln254_unr76_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 14.13 58.56 14.158 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_4_

   PIN memread_edit_dist_g2_ln254_unr76_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 57.202 58.56 57.23 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_5_

   PIN memread_edit_dist_g2_ln254_unr76_q_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.818 0.0 48.846 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_6_

   PIN memread_edit_dist_g2_ln254_unr76_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 2.866 58.56 2.894 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_7_

   PIN memread_edit_dist_g2_ln254_unr76_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 11.314 58.56 11.342 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_9_

   PIN memread_edit_dist_g2_ln254_unr77_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.346 0.0 39.374 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_0_

   PIN memread_edit_dist_g2_ln254_unr77_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.722 0.0 52.75 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_10_

   PIN memread_edit_dist_g2_ln254_unr77_q_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.314 0.0 43.342 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_11_

   PIN memread_edit_dist_g2_ln254_unr77_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.682 0.0 29.71 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_1_

   PIN memread_edit_dist_g2_ln254_unr77_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.202 0.0 41.23 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_2_

   PIN memread_edit_dist_g2_ln254_unr77_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.378 0.0 43.406 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_3_

   PIN memread_edit_dist_g2_ln254_unr77_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.322 0.0 38.35 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_4_

   PIN memread_edit_dist_g2_ln254_unr77_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.746 0.0 29.774 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_5_

   PIN memread_edit_dist_g2_ln254_unr77_q_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.506 0.0 35.534 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_6_

   PIN memread_edit_dist_g2_ln254_unr77_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.89 0.0 43.918 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_7_

   PIN memread_edit_dist_g2_ln254_unr77_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.258 0.0 46.286 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_8_

   PIN memread_edit_dist_g2_ln254_unr77_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 11.122 58.56 11.15 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_9_

   PIN mux_g_ln251_z_911__4472811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.33 0.163 41.358 ;
      END
   END mux_g_ln251_z_911__4472811

   PIN mux_g_ln251_z_923__4472819
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.738 0.163 26.766 ;
      END
   END mux_g_ln251_z_923__4472819

   PIN mux_g_ln251_z_935__4472827
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.186 0.163 11.214 ;
      END
   END mux_g_ln251_z_935__4472827

   PIN mux_g_ln477_q_823_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 39.346 58.56 39.374 ;
      END
   END mux_g_ln477_q_823_

   PIN mux_g_ln477_q_931_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.082 0.0 44.11 0.163 ;
      END
   END mux_g_ln477_q_931_

   PIN n_1796
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 42.674 58.56 42.702 ;
      END
   END n_1796

   PIN n_1809
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 5.746 58.56 5.774 ;
      END
   END n_1809

   PIN n_2052
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 28.594 58.56 28.622 ;
      END
   END n_2052

   PIN n_2059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 14.194 58.56 14.222 ;
      END
   END n_2059

   PIN n_2093
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.69 0.0 56.718 0.163 ;
      END
   END n_2093

   PIN n_2122
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 19.826 58.56 19.854 ;
      END
   END n_2122

   PIN n_21658
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.442 0.163 11.47 ;
      END
   END n_21658

   PIN n_23468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 32.754 58.56 32.782 ;
      END
   END n_23468

   PIN n_23568
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 5.362 58.56 5.39 ;
      END
   END n_23568

   PIN n_23738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 7.922 58.56 7.95 ;
      END
   END n_23738

   PIN n_2401
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 2.93 58.56 2.958 ;
      END
   END n_2401

   PIN n_2442
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.882 0.0 56.91 0.163 ;
      END
   END n_2442

   PIN n_24712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 17.266 58.56 17.294 ;
      END
   END n_24712

   PIN n_25142
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 2.162 58.56 2.19 ;
      END
   END n_25142

   PIN n_25200
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 31.346 58.56 31.374 ;
      END
   END n_25200

   PIN n_2559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 36.21 58.56 36.238 ;
      END
   END n_2559

   PIN n_2653
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 11.506 58.56 11.534 ;
      END
   END n_2653

   PIN n_27360
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.682 0.163 13.71 ;
      END
   END n_27360

   PIN n_29502
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.722 0.082 28.75 ;
      END
   END n_29502

   PIN n_29627
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.482 0.163 42.51 ;
      END
   END n_29627

   PIN n_29628
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.266 0.163 41.294 ;
      END
   END n_29628

   PIN n_29630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.394 0.163 41.422 ;
      END
   END n_29630

   PIN n_29802
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.202 0.163 25.23 ;
      END
   END n_29802

   PIN n_29893
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.842 0.163 25.87 ;
      END
   END n_29893

   PIN n_29895
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.546 0.163 26.574 ;
      END
   END n_29895

   PIN n_30118
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.458 0.163 25.486 ;
      END
   END n_30118

   PIN n_30120
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.61 0.163 26.638 ;
      END
   END n_30120

   PIN n_30316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.554 0.163 45.582 ;
      END
   END n_30316

   PIN n_30339
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.114 0.163 40.142 ;
      END
   END n_30339

   PIN n_30590
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.402 0.163 28.43 ;
      END
   END n_30590

   PIN n_30594
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.338 0.163 28.366 ;
      END
   END n_30594

   PIN n_30671
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.642 0.163 22.67 ;
      END
   END n_30671

   PIN n_30672
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.674 0.163 26.702 ;
      END
   END n_30672

   PIN n_30693
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.05 0.163 24.078 ;
      END
   END n_30693

   PIN n_30772
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.986 0.163 24.014 ;
      END
   END n_30772

   PIN n_30898
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.578 0.163 22.606 ;
      END
   END n_30898

   PIN n_3116
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 14.258 58.56 14.286 ;
      END
   END n_3116

   PIN n_31197
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.186 0.163 75.214 ;
      END
   END n_31197

   PIN n_31199
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.69 0.163 48.718 ;
      END
   END n_31199

   PIN n_31664
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.818 0.163 32.846 ;
      END
   END n_31664

   PIN n_31908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.346 0.163 23.374 ;
      END
   END n_31908

   PIN n_3216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.818 0.0 56.846 0.163 ;
      END
   END n_3216

   PIN n_32226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.114 0.163 72.142 ;
      END
   END n_32226

   PIN n_32312
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.338 0.163 60.366 ;
      END
   END n_32312

   PIN n_32314
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.706 0.163 54.734 ;
      END
   END n_32314

   PIN n_32320
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.618 0.163 69.646 ;
      END
   END n_32320

   PIN n_32321
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.554 0.163 69.582 ;
      END
   END n_32321

   PIN n_32383
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.386 0.163 78.414 ;
      END
   END n_32383

   PIN n_32385
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.994 0.163 43.022 ;
      END
   END n_32385

   PIN n_33478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.882 0.163 16.91 ;
      END
   END n_33478

   PIN n_33638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.522 0.163 57.55 ;
      END
   END n_33638

   PIN n_34651
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.674 0.163 2.702 ;
      END
   END n_34651

   PIN n_34723
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.274 0.082 60.302 ;
      END
   END n_34723

   PIN n_35137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.826 0.163 19.854 ;
      END
   END n_35137

   PIN n_35948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.762 0.163 51.79 ;
      END
   END n_35948

   PIN n_35972
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 74.738 0.163 74.766 ;
      END
   END n_35972

   PIN n_35982
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.69 0.163 48.718 ;
      END
   END n_35982

   PIN n_36120
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.738 0.163 74.766 ;
      END
   END n_36120

   PIN n_36223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 68.722 58.56 68.75 ;
      END
   END n_36223

   PIN n_36620
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.458 0.163 57.486 ;
      END
   END n_36620

   PIN n_36773
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.802 0.163 74.83 ;
      END
   END n_36773

   PIN n_36798
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.506 0.163 35.534 ;
      END
   END n_36798

   PIN n_36805
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.754 0.163 48.782 ;
      END
   END n_36805

   PIN n_36870
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.41 0.163 31.438 ;
      END
   END n_36870

   PIN n_39212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.09 79.837 15.118 80.0 ;
      END
   END n_39212

   PIN n_39292
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.178 0.163 72.206 ;
      END
   END n_39292

   PIN n_39330
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.906 0.163 65.934 ;
      END
   END n_39330

   PIN n_46010
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.986 0.163 8.014 ;
      END
   END n_46010

   PIN n_46011
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.554 0.163 5.582 ;
      END
   END n_46011

   PIN n_49326
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.058 0.163 11.086 ;
      END
   END n_49326

   PIN n_51070
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.162 0.163 66.19 ;
      END
   END n_51070

   PIN n_51313
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.578 0.163 38.606 ;
      END
   END n_51313

   PIN n_51468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.226 0.163 66.254 ;
      END
   END n_51468

   PIN n_52148
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.066 0.163 14.094 ;
      END
   END n_52148

   PIN n_57659
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.466 0.163 60.494 ;
      END
   END n_57659

   PIN n_57660
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.666 0.163 63.694 ;
      END
   END n_57660

   PIN n_58140
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.402 0.163 60.43 ;
      END
   END n_58140

   PIN n_58801
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.13 0.163 14.158 ;
      END
   END n_58801

   PIN n_60533
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.618 0.163 5.646 ;
      END
   END n_60533

   PIN n_61491
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.034 0.163 66.062 ;
      END
   END n_61491

   PIN n_61495
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.922 0.163 39.95 ;
      END
   END n_61495

   PIN n_61496
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.186 0.163 43.214 ;
      END
   END n_61496

   PIN n_62362
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.53 0.163 60.558 ;
      END
   END n_62362

   PIN n_62363
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.898 0.163 62.926 ;
      END
   END n_62363

   PIN n_64805
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.946 0.163 16.974 ;
      END
   END n_64805

   PIN n_65187
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.386 0.0 38.414 0.163 ;
      END
   END n_65187

   PIN n_65196
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 2.674 0.163 2.702 ;
      END
   END n_65196

   PIN n_67247
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.322 0.163 14.35 ;
      END
   END n_67247

   PIN n_8305
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.746 0.163 13.774 ;
      END
   END n_8305

   PIN n_8307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.122 0.163 11.15 ;
      END
   END n_8307

   PIN ternarymux_ln49_0_unr72_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.242 0.163 72.27 ;
      END
   END ternarymux_ln49_0_unr72_z_2_

   PIN ternarymux_ln49_0_unr72_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.306 0.163 72.334 ;
      END
   END ternarymux_ln49_0_unr72_z_3_

   PIN ternarymux_ln49_0_unr76_z_10__4331222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.018 0.163 60.046 ;
      END
   END ternarymux_ln49_0_unr76_z_10__4331222

   PIN ternarymux_ln49_0_unr76_z_8__4331230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.65 0.163 57.678 ;
      END
   END ternarymux_ln49_0_unr76_z_8__4331230

   PIN ternarymux_ln49_0_unr78_z_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.738 0.163 2.766 ;
      END
   END ternarymux_ln49_0_unr78_z_0_

   PIN ternarymux_ln49_0_unr78_z_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.682 0.163 5.71 ;
      END
   END ternarymux_ln49_0_unr78_z_1_

   PIN ternarymux_ln49_0_unr78_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.722 0.163 4.75 ;
      END
   END ternarymux_ln49_0_unr78_z_2_

   PIN ternarymux_ln49_0_unr78_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.05 0.163 8.078 ;
      END
   END ternarymux_ln49_0_unr78_z_3_

   PIN ternarymux_ln49_0_unr78_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.37 0.163 8.398 ;
      END
   END ternarymux_ln49_0_unr78_z_4_

   PIN ternarymux_ln49_0_unr78_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.306 0.163 8.334 ;
      END
   END ternarymux_ln49_0_unr78_z_5_

   PIN ternarymux_ln49_0_unr78_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.21 0.163 20.238 ;
      END
   END ternarymux_ln49_0_unr78_z_6_

   PIN ternarymux_ln49_0_unr78_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.506 0.163 11.534 ;
      END
   END ternarymux_ln49_0_unr78_z_7_

   PIN ternarymux_ln49_0_unr78_z_8__4331262
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.57 0.163 11.598 ;
      END
   END ternarymux_ln49_0_unr78_z_8__4331262

   PIN ternarymux_ln49_0_unr78_z_9__4331258
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.01 0.163 17.038 ;
      END
   END ternarymux_ln49_0_unr78_z_9__4331258

   PIN ternarymux_ln49_5_unr72_z_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.026 0.163 63.054 ;
      END
   END ternarymux_ln49_5_unr72_z_0_

   PIN ternarymux_ln49_6_unr75_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.65 0.163 65.678 ;
      END
   END ternarymux_ln49_6_unr75_z_2_

   PIN ternarymux_ln49_6_unr78_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.25 0.163 11.278 ;
      END
   END ternarymux_ln49_6_unr78_z_12_

   PIN ternarymux_ln49_unr77_z_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.706 0.163 22.734 ;
      END
   END ternarymux_ln49_unr77_z_8_

   PIN FE_OCPN56260_ctrlor_ln251_z_0__4471604_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 7.986 58.56 8.014 ;
      END
   END FE_OCPN56260_ctrlor_ln251_z_0__4471604_bar

   PIN FE_OCPN57864_n_93
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 77.554 58.56 77.582 ;
      END
   END FE_OCPN57864_n_93

   PIN FE_OCPN62021_FE_OFN50813_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 26.546 58.56 26.574 ;
      END
   END FE_OCPN62021_FE_OFN50813_n_67216

   PIN FE_OCPN62025_FE_OFN50813_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 14.45 58.56 14.478 ;
      END
   END FE_OCPN62025_FE_OFN50813_n_67216

   PIN FE_OCPN62349_n_65199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 42.802 58.56 42.83 ;
      END
   END FE_OCPN62349_n_65199

   PIN FE_OCPN62379_FE_OFN47982_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 14.386 58.56 14.414 ;
      END
   END FE_OCPN62379_FE_OFN47982_n_23035

   PIN FE_OCPN62552_FE_OFN47982_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.442 0.0 35.47 0.163 ;
      END
   END FE_OCPN62552_FE_OFN47982_n_23035

   PIN FE_OCPN62858_n_33487_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 8.37 58.56 8.398 ;
      END
   END FE_OCPN62858_n_33487_bar

   PIN FE_OCPN76859_FE_OFN48337_n_31639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.682 79.837 29.71 80.0 ;
      END
   END FE_OCPN76859_FE_OFN48337_n_31639

   PIN FE_OCPN76904_n_58046
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 45.746 58.56 45.774 ;
      END
   END FE_OCPN76904_n_58046

   PIN FE_OCPN77874_FE_OFN48363_n_31641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.802 79.837 2.83 80.0 ;
      END
   END FE_OCPN77874_FE_OFN48363_n_31641

   PIN FE_OFN28531_n_36394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.322 79.837 38.35 80.0 ;
      END
   END FE_OFN28531_n_36394

   PIN FE_OFN28589_n_36353
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.338 79.837 44.366 80.0 ;
      END
   END FE_OFN28589_n_36353

   PIN FE_OFN28736_n_59342
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 13.874 58.56 13.902 ;
      END
   END FE_OFN28736_n_59342

   PIN FE_OFN30021_n_36839
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 72.626 58.56 72.654 ;
      END
   END FE_OFN30021_n_36839

   PIN FE_OFN30124_n_36029
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.234 0.163 37.262 ;
      END
   END FE_OFN30124_n_36029

   PIN FE_OFN30126_n_36012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.978 0.163 37.006 ;
      END
   END FE_OFN30126_n_36012

   PIN FE_OFN30134_n_35994
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.002 0.163 38.03 ;
      END
   END FE_OFN30134_n_35994

   PIN FE_OFN30141_n_34781
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.478 20.274 58.56 20.302 ;
      END
   END FE_OFN30141_n_34781

   PIN FE_OFN30157_n_36428
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.474 0.0 7.502 0.163 ;
      END
   END FE_OFN30157_n_36428

   PIN FE_OFN30217_n_36501
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 7.73 58.56 7.758 ;
      END
   END FE_OFN30217_n_36501

   PIN FE_OFN30294_n_36448
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.266 0.0 41.294 0.163 ;
      END
   END FE_OFN30294_n_36448

   PIN FE_OFN30298_n_36432
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.826 0.0 51.854 0.163 ;
      END
   END FE_OFN30298_n_36432

   PIN FE_OFN30300_n_36379
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 49.65 0.0 49.678 0.163 ;
      END
   END FE_OFN30300_n_36379

   PIN FE_OFN30384_n_34771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 48.69 58.56 48.718 ;
      END
   END FE_OFN30384_n_34771

   PIN FE_OFN30485_n_34770
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 51.442 58.56 51.47 ;
      END
   END FE_OFN30485_n_34770

   PIN FE_OFN30528_n_36408
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 11.314 58.56 11.342 ;
      END
   END FE_OFN30528_n_36408

   PIN FE_OFN30575_n_36929
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.562 0.0 32.59 0.163 ;
      END
   END FE_OFN30575_n_36929

   PIN FE_OFN30593_n_36874
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 14.002 58.56 14.03 ;
      END
   END FE_OFN30593_n_36874

   PIN FE_OFN30767_n_34754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.478 20.722 58.56 20.75 ;
      END
   END FE_OFN30767_n_34754

   PIN FE_OFN30784_n_34754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.258 79.837 38.286 80.0 ;
      END
   END FE_OFN30784_n_34754

   PIN FE_OFN30785_n_34754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.478 4.722 58.56 4.75 ;
      END
   END FE_OFN30785_n_34754

   PIN FE_OFN30819_n_36961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.802 0.0 26.83 0.163 ;
      END
   END FE_OFN30819_n_36961

   PIN FE_OFN30851_n_36114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.858 0.0 15.886 0.163 ;
      END
   END FE_OFN30851_n_36114

   PIN FE_OFN30860_n_34779
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 16.946 58.56 16.974 ;
      END
   END FE_OFN30860_n_34779

   PIN FE_OFN32392_n_51426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 17.65 58.56 17.678 ;
      END
   END FE_OFN32392_n_51426

   PIN FE_OFN32394_n_46215
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.642 58.56 22.67 ;
      END
   END FE_OFN32394_n_46215

   PIN FE_OFN32422_n_62230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.074 0.082 41.102 ;
      END
   END FE_OFN32422_n_62230

   PIN FE_OFN32426_g2_bridge200_rtl_ce_en_3754908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.738 0.163 42.766 ;
      END
   END FE_OFN32426_g2_bridge200_rtl_ce_en_3754908

   PIN FE_OFN34918_n_51730
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 55.026 58.56 55.054 ;
      END
   END FE_OFN34918_n_51730

   PIN FE_OFN34931_n_51721
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 38.002 58.56 38.03 ;
      END
   END FE_OFN34931_n_51721

   PIN FE_OFN34933_memwrite_edit_dist_g2_ln280_unr78_en_0__4469092
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.146 0.163 20.174 ;
      END
   END FE_OFN34933_memwrite_edit_dist_g2_ln280_unr78_en_0__4469092

   PIN FE_OFN35565_n_48865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 39.282 58.56 39.31 ;
      END
   END FE_OFN35565_n_48865

   PIN FE_OFN41927_n_230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.73 79.837 55.758 80.0 ;
      END
   END FE_OFN41927_n_230

   PIN FE_OFN42046_n_232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 5.682 58.56 5.71 ;
      END
   END FE_OFN42046_n_232

   PIN FE_OFN42135_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.002 0.0 54.03 0.163 ;
      END
   END FE_OFN42135_n_222

   PIN FE_OFN42586_n_29
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.818 0.0 48.846 0.163 ;
      END
   END FE_OFN42586_n_29

   PIN FE_OFN42590_n_29
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.106 0.0 21.134 0.163 ;
      END
   END FE_OFN42590_n_29

   PIN FE_OFN42976_n_35330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 54.258 58.56 54.286 ;
      END
   END FE_OFN42976_n_35330

   PIN FE_OFN43000_n_35325
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 52.722 58.56 52.75 ;
      END
   END FE_OFN43000_n_35325

   PIN FE_OFN43003_n_35325
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 55.282 58.56 55.31 ;
      END
   END FE_OFN43003_n_35325

   PIN FE_OFN43167_n_35301
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 33.522 58.56 33.55 ;
      END
   END FE_OFN43167_n_35301

   PIN FE_OFN43216_n_35283
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.434 0.0 56.462 0.163 ;
      END
   END FE_OFN43216_n_35283

   PIN FE_OFN43225_n_35284
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 19.954 58.56 19.982 ;
      END
   END FE_OFN43225_n_35284

   PIN FE_OFN43271_n_35276
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.478 20.146 58.56 20.174 ;
      END
   END FE_OFN43271_n_35276

   PIN FE_OFN43925_mux_g_ln477_q_821_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 55.346 58.56 55.374 ;
      END
   END FE_OFN43925_mux_g_ln477_q_821_

   PIN FE_OFN43998_n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 17.586 58.56 17.614 ;
      END
   END FE_OFN43998_n_35331

   PIN FE_OFN46306_n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 71.922 58.56 71.95 ;
      END
   END FE_OFN46306_n_35331

   PIN FE_OFN47138_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.306 0.0 48.334 0.163 ;
      END
   END FE_OFN47138_n_23039

   PIN FE_OFN47317_n_35285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 42.61 58.56 42.638 ;
      END
   END FE_OFN47317_n_35285

   PIN FE_OFN47849_n_23045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 74.674 58.56 74.702 ;
      END
   END FE_OFN47849_n_23045

   PIN FE_OFN48291_n_31625
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.634 79.837 51.662 80.0 ;
      END
   END FE_OFN48291_n_31625

   PIN FE_OFN48300_n_31625
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.562 79.837 32.59 80.0 ;
      END
   END FE_OFN48300_n_31625

   PIN FE_OFN48307_n_31634
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.538 0.163 71.566 ;
      END
   END FE_OFN48307_n_31634

   PIN FE_OFN48343_n_31639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.314 79.837 3.342 80.0 ;
      END
   END FE_OFN48343_n_31639

   PIN FE_OFN48353_n_31638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.802 79.837 26.83 80.0 ;
      END
   END FE_OFN48353_n_31638

   PIN FE_OFN48358_n_31637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.042 0.163 45.07 ;
      END
   END FE_OFN48358_n_31637

   PIN FE_OFN48629_n_31308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.282 79.837 39.31 80.0 ;
      END
   END FE_OFN48629_n_31308

   PIN FE_OFN48687_n_59052
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.01 79.837 57.038 80.0 ;
      END
   END FE_OFN48687_n_59052

   PIN FE_OFN49699_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 72.562 58.56 72.59 ;
      END
   END FE_OFN49699_n_87

   PIN FE_OFN49700_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 45.874 58.56 45.902 ;
      END
   END FE_OFN49700_n_87

   PIN FE_OFN50548_lt_ln49_6_unr78_z
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.65 0.082 17.678 ;
      END
   END FE_OFN50548_lt_ln49_6_unr78_z

   PIN FE_OFN50882_n_35300
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.714 0.0 41.742 0.163 ;
      END
   END FE_OFN50882_n_35300

   PIN FE_OFN51004_n_23330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 13.938 58.56 13.966 ;
      END
   END FE_OFN51004_n_23330

   PIN FE_OFN53892_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.85 0.0 52.878 0.082 ;
      END
   END FE_OFN53892_n_71

   PIN FE_OFN55363_n_59053
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.618 79.837 29.646 80.0 ;
      END
   END FE_OFN55363_n_59053

   PIN FE_OFN64277_n_57747
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 78.45 58.56 78.478 ;
      END
   END FE_OFN64277_n_57747

   PIN FE_OFN70360_n_36808
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.714 79.837 49.742 80.0 ;
      END
   END FE_OFN70360_n_36808

   PIN FE_OFN70362_n_36328
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.274 0.163 60.302 ;
      END
   END FE_OFN70362_n_36328

   PIN FE_OFN71104_memwrite_edit_dist_g2_ln280_unr73_en_0__4469519
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 54.45 58.56 54.478 ;
      END
   END FE_OFN71104_memwrite_edit_dist_g2_ln280_unr73_en_0__4469519

   PIN FE_OFN71829_n_53368
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 74.674 58.56 74.702 ;
      END
   END FE_OFN71829_n_53368

   PIN FE_OFN73300_n_57
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.978 0.0 53.006 0.163 ;
      END
   END FE_OFN73300_n_57

   PIN FE_OFN73345_n_41
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 68.786 58.56 68.814 ;
      END
   END FE_OFN73345_n_41

   PIN FE_OFN74070_n_59125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.498 79.837 32.526 80.0 ;
      END
   END FE_OFN74070_n_59125

   PIN FE_OFN74248_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 32.818 58.56 32.846 ;
      END
   END FE_OFN74248_n_223

   PIN FE_OFN74309_n_61
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.842 0.0 49.87 0.163 ;
      END
   END FE_OFN74309_n_61

   PIN FE_OFN74356_n_86
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.738 79.837 26.766 80.0 ;
      END
   END FE_OFN74356_n_86

   PIN FE_OFN74575_n_93
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 57.01 79.837 57.038 80.0 ;
      END
   END FE_OFN74575_n_93

   PIN FE_OFN74579_n_79
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.37 79.837 56.398 80.0 ;
      END
   END FE_OFN74579_n_79

   PIN FE_OFN74596_n_856
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.938 0.0 45.966 0.163 ;
      END
   END FE_OFN74596_n_856

   PIN FE_OFN74836_n_34785
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 73.842 58.56 73.87 ;
      END
   END FE_OFN74836_n_34785

   PIN FE_OFN75116_n_34732
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 42.482 58.56 42.51 ;
      END
   END FE_OFN75116_n_34732

   PIN FE_OFN75232_n_35287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 45.682 58.56 45.71 ;
      END
   END FE_OFN75232_n_35287

   PIN FE_OFN75274_n_35301
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.394 79.837 49.422 80.0 ;
      END
   END FE_OFN75274_n_35301

   PIN FE_OFN83829_n_36361
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.026 79.837 39.054 80.0 ;
      END
   END FE_OFN83829_n_36361

   PIN FE_OFN84036_n_7936
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 8.562 58.56 8.59 ;
      END
   END FE_OFN84036_n_7936

   PIN FE_OFN85095_n_30
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.442 79.837 35.47 80.0 ;
      END
   END FE_OFN85095_n_30

   PIN FE_OFN85116_n_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.626 0.0 56.654 0.163 ;
      END
   END FE_OFN85116_n_15

   PIN FE_OFN85912_ternarymux_ln49_0_unr75_z_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.602 0.163 63.63 ;
      END
   END FE_OFN85912_ternarymux_ln49_0_unr75_z_1_

   PIN FE_OFN86076_n_59125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.21 79.837 12.238 80.0 ;
      END
   END FE_OFN86076_n_59125

   PIN FE_OFN86112_mux_g_ln251_z_933__4472823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 10.482 58.56 10.51 ;
      END
   END FE_OFN86112_mux_g_ln251_z_933__4472823

   PIN FE_OFN86557_n_36439
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.498 0.0 32.526 0.163 ;
      END
   END FE_OFN86557_n_36439

   PIN FE_OFN86620_n_35995
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.018 0.0 44.046 0.163 ;
      END
   END FE_OFN86620_n_35995

   PIN FE_OFN86638_n_36832
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.378 0.0 35.406 0.163 ;
      END
   END FE_OFN86638_n_36832

   PIN FE_OFN86665_n_36390
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.898 58.56 22.926 ;
      END
   END FE_OFN86665_n_36390

   PIN FE_OFN86720_n_36698
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 47.602 58.56 47.63 ;
      END
   END FE_OFN86720_n_36698

   PIN FE_OFN86741_n_37010
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 25.65 58.56 25.678 ;
      END
   END FE_OFN86741_n_37010

   PIN FE_OFN86745_n_36401
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 42.866 58.56 42.894 ;
      END
   END FE_OFN86745_n_36401

   PIN FE_OFN86746_n_36399
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.178 0.0 48.206 0.163 ;
      END
   END FE_OFN86746_n_36399

   PIN FE_OFN86876_n_37029
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 2.674 58.56 2.702 ;
      END
   END FE_OFN86876_n_37029

   PIN FE_OFN86890_n_37046
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 41.906 58.56 41.934 ;
      END
   END FE_OFN86890_n_37046

   PIN FE_OFN86897_n_36447
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.834 58.56 22.862 ;
      END
   END FE_OFN86897_n_36447

   PIN FE_OFN87024_n_34784
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 35.442 58.56 35.47 ;
      END
   END FE_OFN87024_n_34784

   PIN FE_OFN88035_mux_g_ln477_q_848_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 17.01 58.56 17.038 ;
      END
   END FE_OFN88035_mux_g_ln477_q_848_

   PIN FE_OFN88305_n_65239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 69.362 58.56 69.39 ;
      END
   END FE_OFN88305_n_65239

   PIN FE_OFN88312_n_65240
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 42.738 58.56 42.766 ;
      END
   END FE_OFN88312_n_65240

   PIN FE_OFN88350_n_26962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.978 0.163 69.006 ;
      END
   END FE_OFN88350_n_26962

   PIN FE_OFN89020_n_31626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.778 0.163 65.806 ;
      END
   END FE_OFN89020_n_31626

   PIN FE_OFN89196_FE_OCPN63783_FE_OFN48830_n_31626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.098 79.837 18.126 80.0 ;
      END
   END FE_OFN89196_FE_OCPN63783_FE_OFN48830_n_31626

   PIN FE_OFN90979_n_22947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 14.322 58.56 14.35 ;
      END
   END FE_OFN90979_n_22947

   PIN FE_OFN95872_n_58716
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.77 58.56 22.798 ;
      END
   END FE_OFN95872_n_58716

   PIN FE_OFN98488_n_35997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 34.354 58.56 34.382 ;
      END
   END FE_OFN98488_n_35997

   PIN FE_OFN98505_n_36246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.042 0.0 53.07 0.163 ;
      END
   END FE_OFN98505_n_36246

   PIN FE_OFN98507_n_36073
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.002 58.56 22.03 ;
      END
   END FE_OFN98507_n_36073

   PIN FE_OFN98899_n_35297
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.066 79.837 54.094 80.0 ;
      END
   END FE_OFN98899_n_35297

   PIN FE_RN_2506_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.29 0.163 50.318 ;
      END
   END FE_RN_2506_0

   PIN FE_RN_3497_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.842 0.163 65.87 ;
      END
   END FE_RN_3497_0

   PIN FE_RN_4443_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.394 0.163 57.422 ;
      END
   END FE_RN_4443_0

   PIN FE_RN_4457_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 43.058 0.163 43.086 ;
      END
   END FE_RN_4457_0

   PIN a_in_104_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.194 0.163 14.222 ;
      END
   END a_in_104_3

   PIN a_in_71_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.594 0.163 28.622 ;
      END
   END a_in_71_3

   PIN a_in_73_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.474 0.163 31.502 ;
      END
   END a_in_73_3

   PIN a_in_78_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.706 0.163 14.734 ;
      END
   END a_in_78_0

   PIN a_in_81_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 32.626 0.163 32.654 ;
      END
   END a_in_81_2

   PIN a_in_87_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.714 0.163 25.742 ;
      END
   END a_in_87_3

   PIN add_85528_72_n_1794471
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.146 0.163 36.174 ;
      END
   END add_85528_72_n_1794471

   PIN add_85528_72_n_4327661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 37.17 0.163 37.198 ;
      END
   END add_85528_72_n_4327661

   PIN add_ln174_1_unr75_z_8__2227682
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.498 0.163 48.526 ;
      END
   END add_ln174_1_unr75_z_8__2227682

   PIN b_in_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.778 79.837 49.806 80.0 ;
      END
   END b_in_2_3

   PIN g2_q69_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.602 0.163 31.63 ;
      END
   END g2_q69_10_

   PIN g2_q69_1__4327571
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.218 0.163 31.246 ;
      END
   END g2_q69_1__4327571

   PIN g2_q69_2__4327573
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 19.89 0.163 19.918 ;
      END
   END g2_q69_2__4327573

   PIN g2_q69_3__4327574
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.162 0.163 34.19 ;
      END
   END g2_q69_3__4327574

   PIN g2_q69_5__4327578
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.538 0.163 31.566 ;
      END
   END g2_q69_5__4327578

   PIN g2_q69_7__4327567
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 37.234 0.163 37.262 ;
      END
   END g2_q69_7__4327567

   PIN g2_q70_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.922 0.163 7.95 ;
      END
   END g2_q70_10_

   PIN g2_q70_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.506 0.163 51.534 ;
      END
   END g2_q70_11_

   PIN g2_q70_3__4327605
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.85 0.163 36.878 ;
      END
   END g2_q70_3__4327605

   PIN g2_q70_5__4327609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.858 0.163 39.886 ;
      END
   END g2_q70_5__4327609

   PIN g2_q70_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.794 0.163 39.822 ;
      END
   END g2_q70_8_

   PIN g2_q71_4__4327638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.754 0.163 48.782 ;
      END
   END g2_q71_4__4327638

   PIN g2_q71_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.618 0.163 45.646 ;
      END
   END g2_q71_8_

   PIN g2_q72_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.482 0.163 10.51 ;
      END
   END g2_q72_10_

   PIN g2_q72_2__4327665
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.082 0.163 36.11 ;
      END
   END g2_q72_2__4327665

   PIN g2_q72_3__4327666
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.722 0.163 36.75 ;
      END
   END g2_q72_3__4327666

   PIN g2_q72_5__4327670
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.746 0.163 29.774 ;
      END
   END g2_q72_5__4327670

   PIN g2_q72_6__4327658
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.114 0.163 40.142 ;
      END
   END g2_q72_6__4327658

   PIN g2_q72_7__4327659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 29.682 0.163 29.71 ;
      END
   END g2_q72_7__4327659

   PIN g2_q73_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 42.866 0.163 42.894 ;
      END
   END g2_q73_11_

   PIN g2_q73_3__4327696
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.45 0.163 78.478 ;
      END
   END g2_q73_3__4327696

   PIN g2_q73_5__4327700
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.378 0.163 51.406 ;
      END
   END g2_q73_5__4327700

   PIN g2_q73_6__4327688
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.05 0.163 40.078 ;
      END
   END g2_q73_6__4327688

   PIN g2_q73_7__4327689
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.21 0.163 60.238 ;
      END
   END g2_q73_7__4327689

   PIN g2_q74_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.122 0.163 75.15 ;
      END
   END g2_q74_11_

   PIN g2_q74_4__4327730
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 75.122 0.163 75.15 ;
      END
   END g2_q74_4__4327730

   PIN g2_q74_5__4327731
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.946 0.163 72.974 ;
      END
   END g2_q74_5__4327731

   PIN g2_q77_2__4327816
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.818 79.837 32.846 80.0 ;
      END
   END g2_q77_2__4327816

   PIN gt_93958_62_n_148_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.394 0.163 57.422 ;
      END
   END gt_93958_62_n_148_bar

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 49.522 0.0 49.55 0.082 ;
      END
   END ispd_clk

   PIN memread_edit_dist_a_ln268_unr124_a_9__4329837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 31.282 58.56 31.31 ;
      END
   END memread_edit_dist_a_ln268_unr124_a_9__4329837

   PIN memread_edit_dist_g2_ln254_unr66_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.29 0.163 34.318 ;
      END
   END memread_edit_dist_g2_ln254_unr66_q_11_

   PIN memread_edit_dist_g2_ln254_unr67_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.954 0.0 43.982 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr67_q_6_

   PIN memread_edit_dist_g2_ln254_unr68_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.746 0.163 45.774 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_0_

   PIN memread_edit_dist_g2_ln254_unr68_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.122 0.163 43.15 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_4_

   PIN memread_edit_dist_g2_ln254_unr68_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.882 0.163 48.91 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_7_

   PIN memread_edit_dist_g2_ln254_unr69_q_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 35.442 0.163 35.47 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_10_

   PIN memread_edit_dist_g2_ln254_unr69_q_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.242 0.0 48.27 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_3_

   PIN memread_edit_dist_g2_ln254_unr69_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.898 0.0 46.926 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_6_

   PIN memread_edit_dist_g2_ln254_unr69_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.722 0.0 52.75 0.163 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_7_

   PIN memread_edit_dist_g2_ln254_unr70_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 19.506 58.56 19.534 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_11_

   PIN memread_edit_dist_g2_ln254_unr70_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.082 0.163 20.11 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_8_

   PIN memwrite_edit_dist_g2_ln280_unr75_en_0__4469773
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.914 0.163 68.942 ;
      END
   END memwrite_edit_dist_g2_ln280_unr75_en_0__4469773

   PIN memwrite_edit_dist_g2_ln280_unr76_en_0__4469257
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.338 0.163 44.366 ;
      END
   END memwrite_edit_dist_g2_ln280_unr76_en_0__4469257

   PIN mux_g_ln477_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.586 79.837 49.614 80.0 ;
      END
   END mux_g_ln477_q_11_

   PIN mux_g_ln477_q_520_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 38.578 58.56 38.606 ;
      END
   END mux_g_ln477_q_520_

   PIN mux_g_ln477_q_799_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 34.226 58.56 34.254 ;
      END
   END mux_g_ln477_q_799_

   PIN mux_g_ln477_q_803_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 19.762 58.56 19.79 ;
      END
   END mux_g_ln477_q_803_

   PIN mux_g_ln477_q_806_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.106 0.0 53.134 0.163 ;
      END
   END mux_g_ln477_q_806_

   PIN mux_g_ln477_q_810_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 11.25 58.56 11.278 ;
      END
   END mux_g_ln477_q_810_

   PIN mux_g_ln477_q_811_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 19.698 58.56 19.726 ;
      END
   END mux_g_ln477_q_811_

   PIN mux_g_ln477_q_814_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 8.306 58.56 8.334 ;
      END
   END mux_g_ln477_q_814_

   PIN mux_g_ln477_q_815_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 19.634 58.56 19.662 ;
      END
   END mux_g_ln477_q_815_

   PIN mux_g_ln477_q_816_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.858 0.0 55.886 0.163 ;
      END
   END mux_g_ln477_q_816_

   PIN mux_g_ln477_q_818_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 51.506 58.56 51.534 ;
      END
   END mux_g_ln477_q_818_

   PIN mux_g_ln477_q_820_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.914 0.0 52.942 0.163 ;
      END
   END mux_g_ln477_q_820_

   PIN mux_g_ln477_q_827_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 8.242 58.56 8.27 ;
      END
   END mux_g_ln477_q_827_

   PIN mux_g_ln477_q_831_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 49.778 0.0 49.806 0.163 ;
      END
   END mux_g_ln477_q_831_

   PIN mux_g_ln477_q_834_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 8.178 58.56 8.206 ;
      END
   END mux_g_ln477_q_834_

   PIN mux_g_ln477_q_835_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 36.146 58.56 36.174 ;
      END
   END mux_g_ln477_q_835_

   PIN mux_g_ln477_q_836_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 26.482 58.56 26.51 ;
      END
   END mux_g_ln477_q_836_

   PIN mux_g_ln477_q_841_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.818 0.0 56.846 0.163 ;
      END
   END mux_g_ln477_q_841_

   PIN mux_g_ln477_q_846_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 29.682 58.56 29.71 ;
      END
   END mux_g_ln477_q_846_

   PIN mux_g_ln477_q_851_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 5.618 58.56 5.646 ;
      END
   END mux_g_ln477_q_851_

   PIN n_21259
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 41.842 58.56 41.87 ;
      END
   END n_21259

   PIN n_21278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 38.77 58.56 38.798 ;
      END
   END n_21278

   PIN n_21287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 66.802 58.56 66.83 ;
      END
   END n_21287

   PIN n_23142
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 30.322 58.56 30.35 ;
      END
   END n_23142

   PIN n_23298
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.802 0.163 34.83 ;
      END
   END n_23298

   PIN n_23337
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.242 0.163 32.27 ;
      END
   END n_23337

   PIN n_23348
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.258 0.0 30.286 0.163 ;
      END
   END n_23348

   PIN n_26820
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.042 0.163 69.07 ;
      END
   END n_26820

   PIN n_27167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.49 0.163 69.518 ;
      END
   END n_27167

   PIN n_27169
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.09 0.163 63.118 ;
      END
   END n_27169

   PIN n_27172
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.322 0.163 78.35 ;
      END
   END n_27172

   PIN n_27478
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.722 0.082 68.75 ;
      END
   END n_27478

   PIN n_28223
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.97 0.163 65.998 ;
      END
   END n_28223

   PIN n_28405
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.522 0.082 65.55 ;
      END
   END n_28405

   PIN n_28469
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.426 0.163 69.454 ;
      END
   END n_28469

   PIN n_28821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.65 0.0 49.678 0.163 ;
      END
   END n_28821

   PIN n_28879
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.01 0.0 49.038 0.163 ;
      END
   END n_28879

   PIN n_29799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.202 0.163 41.23 ;
      END
   END n_29799

   PIN n_30353
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.234 0.082 45.262 ;
      END
   END n_30353

   PIN n_3063
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.938 0.163 13.966 ;
      END
   END n_3063

   PIN n_30960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.682 0.163 29.71 ;
      END
   END n_30960

   PIN n_30965
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.106 0.163 29.134 ;
      END
   END n_30965

   PIN n_31888
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.354 0.163 50.382 ;
      END
   END n_31888

   PIN n_32070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.93 0.163 34.958 ;
      END
   END n_32070

   PIN n_32511
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.33 0.163 57.358 ;
      END
   END n_32511

   PIN n_33240
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.098 0.163 50.126 ;
      END
   END n_33240

   PIN n_33245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.778 0.163 17.806 ;
      END
   END n_33245

   PIN n_33384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.442 0.163 51.47 ;
      END
   END n_33384

   PIN n_33386
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.322 0.163 54.35 ;
      END
   END n_33386

   PIN n_33467_bar
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 8.114 58.56 8.142 ;
      END
   END n_33467_bar

   PIN n_33556
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.762 0.163 59.79 ;
      END
   END n_33556

   PIN n_33599
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.826 0.163 59.854 ;
      END
   END n_33599

   PIN n_33639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.522 0.163 49.55 ;
      END
   END n_33639

   PIN n_3370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 36.722 58.56 36.75 ;
      END
   END n_3370

   PIN n_34235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.258 0.163 54.286 ;
      END
   END n_34235

   PIN n_34404
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.522 0.082 17.55 ;
      END
   END n_34404

   PIN n_34535
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.578 0.163 62.606 ;
      END
   END n_34535

   PIN n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 16.882 58.56 16.91 ;
      END
   END n_35331

   PIN n_35936
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.85 0.0 52.878 0.163 ;
      END
   END n_35936

   PIN n_35978
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.706 58.56 22.734 ;
      END
   END n_35978

   PIN n_35984
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.154 0.0 55.182 0.163 ;
      END
   END n_35984

   PIN n_36005
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 54.386 58.56 54.414 ;
      END
   END n_36005

   PIN n_36014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 5.554 58.56 5.582 ;
      END
   END n_36014

   PIN n_36015
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 32.242 58.56 32.27 ;
      END
   END n_36015

   PIN n_36035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 16.818 58.56 16.846 ;
      END
   END n_36035

   PIN n_36060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 25.586 58.56 25.614 ;
      END
   END n_36060

   PIN n_36062
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 11.186 58.56 11.214 ;
      END
   END n_36062

   PIN n_36086
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.578 58.56 22.606 ;
      END
   END n_36086

   PIN n_36113
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.026 0.0 23.054 0.163 ;
      END
   END n_36113

   PIN n_36221
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.778 0.0 49.806 0.163 ;
      END
   END n_36221

   PIN n_36250
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 16.882 58.56 16.91 ;
      END
   END n_36250

   PIN n_36339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 8.434 58.56 8.462 ;
      END
   END n_36339

   PIN n_36355
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.834 79.837 30.862 80.0 ;
      END
   END n_36355

   PIN n_36486
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.714 0.0 49.742 0.163 ;
      END
   END n_36486

   PIN n_36520
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 5.746 58.56 5.774 ;
      END
   END n_36520

   PIN n_36547
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.25 0.0 3.278 0.163 ;
      END
   END n_36547

   PIN n_36563
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 37.042 58.56 37.07 ;
      END
   END n_36563

   PIN n_36622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 11.058 58.56 11.086 ;
      END
   END n_36622

   PIN n_36733
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 2.674 58.56 2.702 ;
      END
   END n_36733

   PIN n_36748
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 13.682 58.56 13.71 ;
      END
   END n_36748

   PIN n_36785
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 36.082 58.56 36.11 ;
      END
   END n_36785

   PIN n_36787
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 19.57 58.56 19.598 ;
      END
   END n_36787

   PIN n_36803
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.674 0.0 50.702 0.163 ;
      END
   END n_36803

   PIN n_36899
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 22.514 58.56 22.542 ;
      END
   END n_36899

   PIN n_36922
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 16.754 58.56 16.782 ;
      END
   END n_36922

   PIN n_36928
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 42.546 58.56 42.574 ;
      END
   END n_36928

   PIN n_36944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.602 0.0 55.63 0.163 ;
      END
   END n_36944

   PIN n_36948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.962 0.0 54.99 0.163 ;
      END
   END n_36948

   PIN n_36953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 16.69 58.56 16.718 ;
      END
   END n_36953

   PIN n_36965
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 16.626 58.56 16.654 ;
      END
   END n_36965

   PIN n_36980
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.258 0.0 38.286 0.163 ;
      END
   END n_36980

   PIN n_39130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.754 0.163 16.782 ;
      END
   END n_39130

   PIN n_39362
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.922 0.163 7.95 ;
      END
   END n_39362

   PIN n_42401
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.914 0.163 36.942 ;
      END
   END n_42401

   PIN n_43309
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.45 0.082 62.478 ;
      END
   END n_43309

   PIN n_45751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.962 0.163 62.99 ;
      END
   END n_45751

   PIN n_45752
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.562 79.837 24.59 80.0 ;
      END
   END n_45752

   PIN n_46296
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.274 79.837 12.302 80.0 ;
      END
   END n_46296

   PIN n_51091
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 65.522 58.56 65.55 ;
      END
   END n_51091

   PIN n_53413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 46.962 58.56 46.99 ;
      END
   END n_53413

   PIN n_56864
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.322 0.163 62.35 ;
      END
   END n_56864

   PIN n_56944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.402 79.837 52.43 80.0 ;
      END
   END n_56944

   PIN n_57
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.162 0.0 18.19 0.163 ;
      END
   END n_57

   PIN n_57749
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 51.57 58.56 51.598 ;
      END
   END n_57749

   PIN n_57753
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 48.818 58.56 48.846 ;
      END
   END n_57753

   PIN n_58050
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 48.754 58.56 48.782 ;
      END
   END n_58050

   PIN n_58450
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.082 79.837 44.11 80.0 ;
      END
   END n_58450

   PIN n_58539
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.666 79.837 55.694 80.0 ;
      END
   END n_58539

   PIN n_58771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 58.397 42.482 58.56 42.51 ;
      END
   END n_58771

   PIN n_58784
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.442 0.163 19.47 ;
      END
   END n_58784

   PIN n_6033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 28.466 58.56 28.494 ;
      END
   END n_6033

   PIN n_60540
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.314 0.163 11.342 ;
      END
   END n_60540

   PIN n_60542
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.49 0.163 21.518 ;
      END
   END n_60542

   PIN n_60548
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.162 0.163 26.19 ;
      END
   END n_60548

   PIN n_60638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.146 0.163 60.174 ;
      END
   END n_60638

   PIN n_64833
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.874 0.082 45.902 ;
      END
   END n_64833

   PIN n_64835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.514 0.082 54.542 ;
      END
   END n_64835

   PIN n_65250
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 58.397 78.322 58.56 78.35 ;
      END
   END n_65250

   PIN n_66515
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.378 0.163 11.406 ;
      END
   END n_66515

   PIN n_67153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.53 0.163 44.558 ;
      END
   END n_67153

   PIN ternarymux_ln49_0_unr72_z_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.386 0.163 54.414 ;
      END
   END ternarymux_ln49_0_unr72_z_1_

   PIN ternarymux_ln49_0_unr75_z_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.05 0.163 72.078 ;
      END
   END ternarymux_ln49_0_unr75_z_0_

   PIN ternarymux_ln49_0_unr75_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.53 0.163 68.558 ;
      END
   END ternarymux_ln49_0_unr75_z_2_

   PIN ternarymux_ln49_0_unr75_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.922 0.163 71.95 ;
      END
   END ternarymux_ln49_0_unr75_z_3_

   PIN ternarymux_ln49_0_unr75_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.986 0.163 72.014 ;
      END
   END ternarymux_ln49_0_unr75_z_4_

   PIN ternarymux_ln49_0_unr75_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.458 0.163 57.486 ;
      END
   END ternarymux_ln49_0_unr75_z_5_

   PIN ternarymux_ln49_0_unr75_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.194 0.163 54.222 ;
      END
   END ternarymux_ln49_0_unr75_z_6_

   PIN ternarymux_ln49_0_unr75_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.13 0.163 54.158 ;
      END
   END ternarymux_ln49_0_unr75_z_7_

   PIN ternarymux_ln49_0_unr76_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.682 0.163 53.71 ;
      END
   END ternarymux_ln49_0_unr76_z_5_

   PIN ternarymux_ln49_0_unr76_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.77 0.163 54.798 ;
      END
   END ternarymux_ln49_0_unr76_z_6_

   PIN ternarymux_ln49_0_unr76_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.082 0.163 52.11 ;
      END
   END ternarymux_ln49_0_unr76_z_7_

   PIN ternarymux_ln49_0_unr76_z_9__4331226
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.682 0.163 45.71 ;
      END
   END ternarymux_ln49_0_unr76_z_9__4331226

   PIN ternarymux_ln49_6_unr77_z_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.042 0.163 29.07 ;
      END
   END ternarymux_ln49_6_unr77_z_8_

   PIN ternarymux_ln49_8_unr72_z_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.466 0.163 68.494 ;
      END
   END ternarymux_ln49_8_unr72_z_0_

   PIN ternarymux_ln49_8_unr72_z_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.594 0.163 68.622 ;
      END
   END ternarymux_ln49_8_unr72_z_1_

   PIN ternarymux_ln49_8_unr78_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.602 0.163 7.63 ;
      END
   END ternarymux_ln49_8_unr78_z_10_

   PIN ternarymux_ln49_unr75_z_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.362 0.163 69.39 ;
      END
   END ternarymux_ln49_unr75_z_0_

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 58.56 80.0 ;
      LAYER V1 ;
         RECT 0.0 0.0 58.56 80.0 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 58.56 80.0 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 58.56 80.0 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 58.56 80.0 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 58.56 80.0 ;
      LAYER M1 ;
         RECT 0.0 0.0 58.56 80.0 ;
   END
END h1_mgc_edit_dist_a

MACRO h4_mgc_matrix_mult_a
   CLASS BLOCK ;
   FOREIGN h4 ;
   ORIGIN 0 0 ;
   SIZE 158.72 BY 106.24 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN11536_n_140234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.506 0.0 35.534 0.082 ;
      END
   END FE_OFN11536_n_140234

   PIN FE_OFN11537_n_140234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.434 0.0 24.462 0.082 ;
      END
   END FE_OFN11537_n_140234

   PIN FE_OFN13236_n_143479
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.698 0.0 27.726 0.163 ;
      END
   END FE_OFN13236_n_143479

   PIN FE_OFN16095_n_143423
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.546 0.0 66.574 0.163 ;
      END
   END FE_OFN16095_n_143423

   PIN FE_OFN18007_n_143669
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.09 0.163 7.118 ;
      END
   END FE_OFN18007_n_143669

   PIN FE_OFN6242_delay_mul_ln34_unr7_unr3_stage2_stallmux_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.106 0.0 101.134 0.163 ;
      END
   END FE_OFN6242_delay_mul_ln34_unr7_unr3_stage2_stallmux_z_5_

   PIN FE_OFN6244_delay_mul_ln34_unr7_unr3_stage2_stallmux_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.882 0.0 128.91 0.163 ;
      END
   END FE_OFN6244_delay_mul_ln34_unr7_unr3_stage2_stallmux_z_4_

   PIN FE_OFN6343_delay_mul_ln34_unr7_unr1_stage2_stallmux_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.922 0.0 143.95 0.163 ;
      END
   END FE_OFN6343_delay_mul_ln34_unr7_unr1_stage2_stallmux_z_6_

   PIN FE_OFN6345_delay_mul_ln34_unr7_unr1_stage2_stallmux_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.73 0.0 151.758 0.163 ;
      END
   END FE_OFN6345_delay_mul_ln34_unr7_unr1_stage2_stallmux_z_5_

   PIN FE_OFN6357_delay_mul_ln34_unr7_unr1_stage2_stallmux_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.898 0.0 110.926 0.163 ;
      END
   END FE_OFN6357_delay_mul_ln34_unr7_unr1_stage2_stallmux_z_4_

   PIN FE_OFN6470_n_137680
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.626 0.163 64.654 ;
      END
   END FE_OFN6470_n_137680

   PIN FE_OFN6472_delay_mul_ln34_unr7_unr3_stage2_stallmux_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.546 0.0 58.574 0.163 ;
      END
   END FE_OFN6472_delay_mul_ln34_unr7_unr3_stage2_stallmux_z_2_

   PIN FE_OFN6474_delay_mul_ln34_unr7_unr3_stage2_stallmux_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.61 0.0 146.638 0.163 ;
      END
   END FE_OFN6474_delay_mul_ln34_unr7_unr3_stage2_stallmux_z_3_

   PIN FE_OFN6561_n_120781
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.13 0.0 70.158 0.163 ;
      END
   END FE_OFN6561_n_120781

   PIN FE_OFN7002_n_140202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.082 0.163 4.11 ;
      END
   END FE_OFN7002_n_140202

   PIN FE_OFN8439_n_27832
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 26.162 0.163 26.19 ;
      END
   END FE_OFN8439_n_27832

   PIN FE_OFN8442_n_6523
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.65 0.0 17.678 0.163 ;
      END
   END FE_OFN8442_n_6523

   PIN FE_OFN8633_n_31042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.042 106.077 5.07 106.24 ;
      END
   END FE_OFN8633_n_31042

   PIN FE_OFN8641_n_29615
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.194 0.163 102.222 ;
      END
   END FE_OFN8641_n_29615

   PIN FE_OFN8647_n_28444
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 91.506 0.163 91.534 ;
      END
   END FE_OFN8647_n_28444

   PIN FE_OFN8655_n_25409
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 99.122 0.163 99.15 ;
      END
   END FE_OFN8655_n_25409

   PIN delay_mul_ln34_unr7_unr1_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.954 0.0 19.982 0.163 ;
      END
   END delay_mul_ln34_unr7_unr1_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr7_unr1_stage2_stallmux_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.93 0.0 2.958 0.163 ;
      END
   END delay_mul_ln34_unr7_unr1_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr7_unr1_stage2_stallmux_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.578 0.0 134.606 0.163 ;
      END
   END delay_mul_ln34_unr7_unr1_stage2_stallmux_z_3_

   PIN delay_mul_ln34_unr7_unr3_stage2_stallmux_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.042 0.163 61.07 ;
      END
   END delay_mul_ln34_unr7_unr3_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr7_unr3_stage2_stallmux_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.874 0.0 101.902 0.163 ;
      END
   END delay_mul_ln34_unr7_unr3_stage2_stallmux_z_6_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.698 0.0 11.726 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_3_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.082 0.163 20.11 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.802 0.163 18.83 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.306 0.163 72.334 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_10_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.026 0.0 15.054 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.146 0.163 4.174 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 76.146 0.163 76.174 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_9_

   PIN mul_4694_72_n_137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.298 0.0 109.326 0.163 ;
      END
   END mul_4694_72_n_137

   PIN mul_4694_72_n_254
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.738 0.0 50.766 0.163 ;
      END
   END mul_4694_72_n_254

   PIN mul_4694_72_n_295
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.442 0.0 59.47 0.163 ;
      END
   END mul_4694_72_n_295

   PIN mul_4694_72_n_296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.89 0.0 59.918 0.163 ;
      END
   END mul_4694_72_n_296

   PIN mul_4694_72_n_331
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.53 0.0 60.558 0.163 ;
      END
   END mul_4694_72_n_331

   PIN n_112396
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.314 0.0 27.342 0.163 ;
      END
   END n_112396

   PIN n_116308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.442 0.0 19.47 0.163 ;
      END
   END n_116308

   PIN n_116312
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.994 0.0 51.022 0.163 ;
      END
   END n_116312

   PIN n_116493
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.386 0.0 62.414 0.163 ;
      END
   END n_116493

   PIN n_116494
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.322 0.0 62.35 0.163 ;
      END
   END n_116494

   PIN n_116575
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.514 0.0 54.542 0.163 ;
      END
   END n_116575

   PIN n_116621
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.074 0.0 25.102 0.163 ;
      END
   END n_116621

   PIN n_116777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.034 0.0 66.062 0.163 ;
      END
   END n_116777

   PIN n_120549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.466 0.0 36.494 0.163 ;
      END
   END n_120549

   PIN n_120739
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.626 0.0 112.654 0.163 ;
      END
   END n_120739

   PIN n_120779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.874 0.0 69.902 0.163 ;
      END
   END n_120779

   PIN n_120782
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.098 0.0 66.126 0.163 ;
      END
   END n_120782

   PIN n_121450
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.282 0.0 39.31 0.163 ;
      END
   END n_121450

   PIN n_124090
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.802 0.0 66.83 0.163 ;
      END
   END n_124090

   PIN n_137682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.242 0.0 16.27 0.163 ;
      END
   END n_137682

   PIN n_15496
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.594 0.0 4.622 0.163 ;
      END
   END n_15496

   PIN n_16158
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.962 0.0 30.99 0.163 ;
      END
   END n_16158

   PIN n_17902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.474 0.0 31.502 0.163 ;
      END
   END n_17902

   PIN n_18036
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.066 0.163 102.094 ;
      END
   END n_18036

   PIN n_18759
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.002 0.163 94.03 ;
      END
   END n_18759

   PIN n_18760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.682 0.163 93.71 ;
      END
   END n_18760

   PIN n_18766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.258 0.163 102.286 ;
      END
   END n_18766

   PIN n_19998
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.49 0.163 69.518 ;
      END
   END n_19998

   PIN n_21785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.762 0.163 11.79 ;
      END
   END n_21785

   PIN n_22637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 95.218 0.163 95.246 ;
      END
   END n_22637

   PIN n_22638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 95.282 0.163 95.31 ;
      END
   END n_22638

   PIN n_22901
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.41 0.0 7.438 0.163 ;
      END
   END n_22901

   PIN n_26674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.962 0.163 102.99 ;
      END
   END n_26674

   PIN n_27108
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 54.642 0.0 54.67 0.163 ;
      END
   END n_27108

   PIN n_27109
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.642 0.0 54.67 0.163 ;
      END
   END n_27109

   PIN n_27295
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 99.186 0.163 99.214 ;
      END
   END n_27295

   PIN n_27896
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 99.25 0.163 99.278 ;
      END
   END n_27896

   PIN n_28225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.378 0.0 35.406 0.163 ;
      END
   END n_28225

   PIN n_28690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 83.762 0.163 83.79 ;
      END
   END n_28690

   PIN n_28700
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.762 0.0 115.79 0.163 ;
      END
   END n_28700

   PIN n_29119
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 87.666 0.163 87.694 ;
      END
   END n_29119

   PIN n_29550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 103.026 0.163 103.054 ;
      END
   END n_29550

   PIN n_29622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.482 0.0 74.51 0.163 ;
      END
   END n_29622

   PIN n_29623
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.546 0.0 74.574 0.163 ;
      END
   END n_29623

   PIN n_29696
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.01 0.0 73.038 0.163 ;
      END
   END n_29696

   PIN n_29943
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 99.314 0.163 99.342 ;
      END
   END n_29943

   PIN n_30272
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.922 0.163 79.95 ;
      END
   END n_30272

   PIN n_30545
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.106 0.163 61.134 ;
      END
   END n_30545

   PIN n_30553
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.242 0.163 72.27 ;
      END
   END n_30553

   PIN n_30641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.178 0.0 16.206 0.163 ;
      END
   END n_30641

   PIN n_31365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.746 0.163 93.774 ;
      END
   END n_31365

   PIN n_31915
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.482 0.163 42.51 ;
      END
   END n_31915

   PIN n_37096
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.802 0.0 50.83 0.163 ;
      END
   END n_37096

   PIN n_37117
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.29 0.0 58.318 0.163 ;
      END
   END n_37117

   PIN n_37415
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.194 0.0 62.222 0.163 ;
      END
   END n_37415

   PIN n_41861
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.522 0.0 41.55 0.163 ;
      END
   END n_41861

   PIN n_43109
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.154 0.0 39.182 0.163 ;
      END
   END n_43109

   PIN n_43425
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.97 0.0 41.998 0.163 ;
      END
   END n_43425

   PIN n_43426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.218 0.0 39.246 0.163 ;
      END
   END n_43426

   PIN n_4535
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.162 0.163 50.19 ;
      END
   END n_4535

   PIN n_4622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.114 0.0 16.142 0.163 ;
      END
   END n_4622

   PIN n_50299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.994 0.0 43.022 0.163 ;
      END
   END n_50299

   PIN n_50332
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.498 0.0 40.526 0.163 ;
      END
   END n_50332

   PIN n_50333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.17 0.0 37.198 0.163 ;
      END
   END n_50333

   PIN n_50502
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.506 0.0 35.534 0.163 ;
      END
   END n_50502

   PIN n_53705
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.25 0.0 35.278 0.163 ;
      END
   END n_53705

   PIN n_53787
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.858 0.0 23.886 0.163 ;
      END
   END n_53787

   PIN n_5576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.41 0.0 39.438 0.163 ;
      END
   END n_5576

   PIN n_62552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.49 0.0 85.518 0.163 ;
      END
   END n_62552

   PIN n_62941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.554 0.0 77.582 0.163 ;
      END
   END n_62941

   PIN n_63426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.618 0.0 77.646 0.163 ;
      END
   END n_63426

   PIN n_64062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.106 0.0 93.134 0.163 ;
      END
   END n_64062

   PIN n_64537
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.17 0.0 93.198 0.163 ;
      END
   END n_64537

   PIN n_71957
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.138 0.0 97.166 0.163 ;
      END
   END n_71957

   PIN n_97280
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.818 0.0 88.846 0.163 ;
      END
   END n_97280

   PIN FE_OFN11525_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.754 0.0 40.782 0.082 ;
      END
   END FE_OFN11525_n_140234

   PIN FE_OFN11533_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.634 0.0 35.662 0.163 ;
      END
   END FE_OFN11533_n_140234

   PIN FE_OFN12010_n_143453
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.122 0.0 43.15 0.163 ;
      END
   END FE_OFN12010_n_143453

   PIN FE_OFN12011_n_143453
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.09 0.0 39.118 0.163 ;
      END
   END FE_OFN12011_n_143453

   PIN FE_OFN12063_n_143423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.338 0.0 12.366 0.163 ;
      END
   END FE_OFN12063_n_143423

   PIN FE_OFN13199_n_137475
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.41 0.0 31.438 0.163 ;
      END
   END FE_OFN13199_n_137475

   PIN FE_OFN13235_n_143479
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.338 0.0 20.366 0.163 ;
      END
   END FE_OFN13235_n_143479

   PIN FE_OFN13254_n_143369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.506 0.0 19.534 0.082 ;
      END
   END FE_OFN13254_n_143369

   PIN FE_OFN13425_n_41709
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.69 0.0 8.718 0.163 ;
      END
   END FE_OFN13425_n_41709

   PIN FE_OFN13786_n_41960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.778 0.0 9.806 0.163 ;
      END
   END FE_OFN13786_n_41960

   PIN FE_OFN14575_n_41015
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.962 0.0 46.99 0.163 ;
      END
   END FE_OFN14575_n_41015

   PIN FE_OFN15028_n_41964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.53 0.163 28.558 ;
      END
   END FE_OFN15028_n_41964

   PIN FE_OFN17927_n_143370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.29 0.0 42.318 0.163 ;
      END
   END FE_OFN17927_n_143370

   PIN FE_OFN18006_n_143669
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.466 0.0 124.494 0.163 ;
      END
   END FE_OFN18006_n_143669

   PIN FE_OFN18963_n_41993
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.154 0.0 63.182 0.163 ;
      END
   END FE_OFN18963_n_41993

   PIN FE_OFN6236_n_137235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.018 0.0 20.046 0.082 ;
      END
   END FE_OFN6236_n_137235

   PIN FE_OFN6289_delay_mul_ln34_unr7_unr1_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.93 0.0 50.958 0.163 ;
      END
   END FE_OFN6289_delay_mul_ln34_unr7_unr1_stage2_stallmux_z_11_

   PIN FE_OFN6488_n_41961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.21 0.163 4.238 ;
      END
   END FE_OFN6488_n_41961

   PIN FE_OFN6551_n_41963
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.786 0.0 4.814 0.163 ;
      END
   END FE_OFN6551_n_41963

   PIN FE_OFN6628_n_41612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.914 0.0 76.942 0.163 ;
      END
   END FE_OFN6628_n_41612

   PIN FE_OFN6662_n_41611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.442 0.082 3.47 ;
      END
   END FE_OFN6662_n_41611

   PIN FE_OFN6862_n_143629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.802 0.0 50.83 0.163 ;
      END
   END FE_OFN6862_n_143629

   PIN FE_OFN6896_n_143493
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.722 0.0 28.75 0.082 ;
      END
   END FE_OFN6896_n_143493

   PIN FE_OFN8989_n_30545
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.746 106.077 13.774 106.24 ;
      END
   END FE_OFN8989_n_30545

   PIN FE_OFN9645_b_7_3_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.642 0.0 22.67 0.163 ;
      END
   END FE_OFN9645_b_7_3_11

   PIN FE_OFN9659_b_7_3_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.386 0.0 22.414 0.163 ;
      END
   END FE_OFN9659_b_7_3_6

   PIN FE_OFN9662_b_7_3_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.402 0.082 28.43 ;
      END
   END FE_OFN9662_b_7_3_5

   PIN FE_OFN9666_b_7_3_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.57 0.0 19.598 0.163 ;
      END
   END FE_OFN9666_b_7_3_4

   PIN FE_OFN9669_b_7_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.09 0.0 47.118 0.163 ;
      END
   END FE_OFN9669_b_7_3_3

   PIN FE_OFN9672_b_7_3_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.93 0.0 50.958 0.082 ;
      END
   END FE_OFN9672_b_7_3_2

   PIN FE_OFN9675_b_7_3_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.61 0.0 42.638 0.163 ;
      END
   END FE_OFN9675_b_7_3_1

   PIN FE_OFN9677_b_7_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.474 0.0 39.502 0.163 ;
      END
   END FE_OFN9677_b_7_3_0

   PIN FE_OFN9678_b_7_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.274 0.0 12.302 0.163 ;
      END
   END FE_OFN9678_b_7_3_0

   PIN FE_OFN9706_b_7_1_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.346 0.0 39.374 0.163 ;
      END
   END FE_OFN9706_b_7_1_5

   PIN FE_OFN9709_b_7_1_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.466 0.0 12.494 0.163 ;
      END
   END FE_OFN9709_b_7_1_4

   PIN FE_OFN9712_b_7_1_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.882 0.0 16.91 0.163 ;
      END
   END FE_OFN9712_b_7_1_3

   PIN FE_OFN9715_b_7_1_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.666 0.0 31.694 0.163 ;
      END
   END FE_OFN9715_b_7_1_2

   PIN FE_OFN9720_b_7_1_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.218 0.0 39.246 0.163 ;
      END
   END FE_OFN9720_b_7_1_1

   PIN FE_OFN9723_b_7_1_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.914 0.0 4.942 0.163 ;
      END
   END FE_OFN9723_b_7_1_0

   PIN delay_mul_ln34_unr6_unr1_stage2_stallmux_q_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.826 0.163 11.854 ;
      END
   END delay_mul_ln34_unr6_unr1_stage2_stallmux_q_10_

   PIN delay_mul_ln34_unr6_unr1_stage2_stallmux_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.962 0.163 6.99 ;
      END
   END delay_mul_ln34_unr6_unr1_stage2_stallmux_q_11_

   PIN delay_mul_ln34_unr6_unr1_stage2_stallmux_q_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.05 0.0 16.078 0.163 ;
      END
   END delay_mul_ln34_unr6_unr1_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr6_unr1_stage2_stallmux_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.762 0.163 27.79 ;
      END
   END delay_mul_ln34_unr6_unr1_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr6_unr1_stage2_stallmux_q_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.162 0.163 34.19 ;
      END
   END delay_mul_ln34_unr6_unr1_stage2_stallmux_q_9_

   PIN delay_mul_ln34_unr6_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.554 0.0 29.582 0.163 ;
      END
   END delay_mul_ln34_unr6_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr7_unr1_stage2_stallmux_q_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.058 0.0 51.086 0.163 ;
      END
   END delay_mul_ln34_unr7_unr1_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr7_unr1_stage2_stallmux_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.578 0.0 54.606 0.163 ;
      END
   END delay_mul_ln34_unr7_unr1_stage2_stallmux_z_10_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.402 0.163 12.43 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_z_3_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.706 0.163 14.734 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr7_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.602 0.0 31.63 0.163 ;
      END
   END delay_mul_ln34_unr7_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr7_unr8_stage2_stallmux_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.626 0.0 8.654 0.163 ;
      END
   END delay_mul_ln34_unr7_unr8_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr7_unr9_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.778 0.0 17.806 0.163 ;
      END
   END delay_mul_ln34_unr7_unr9_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.026 0.0 47.054 0.163 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_10_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.714 0.0 65.742 0.163 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_11_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.258 0.0 62.286 0.163 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.602 0.0 71.63 0.163 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 0.0 25.614 0.163 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_9_

   PIN delay_mul_ln34_unr8_unr3_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.554 0.163 69.582 ;
      END
   END delay_mul_ln34_unr8_unr3_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr8_unr3_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.986 0.0 32.014 0.163 ;
      END
   END delay_mul_ln34_unr8_unr3_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.002 0.163 102.03 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.378 0.0 3.406 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.25 0.0 3.278 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_z_10_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.786 0.0 4.814 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.114 0.0 8.142 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_z_7_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.69 0.0 8.718 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_z_9_

   PIN delay_mul_ln34_unr8_unr9_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.314 0.0 19.342 0.163 ;
      END
   END delay_mul_ln34_unr8_unr9_stage2_stallmux_q_15_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.882 0.0 8.91 0.082 ;
      END
   END ispd_clk

   PIN mul_4694_72_n_114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.402 0.0 12.43 0.163 ;
      END
   END mul_4694_72_n_114

   PIN mul_4694_72_n_294
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.762 0.0 59.79 0.163 ;
      END
   END mul_4694_72_n_294

   PIN mul_4694_72_n_330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.21 0.0 60.238 0.163 ;
      END
   END mul_4694_72_n_330

   PIN mul_4694_72_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.13 0.0 78.158 0.163 ;
      END
   END mul_4694_72_n_50

   PIN mul_4694_72_n_66
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.066 0.0 78.094 0.163 ;
      END
   END mul_4694_72_n_66

   PIN mul_4694_72_n_793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.866 0.0 50.894 0.163 ;
      END
   END mul_4694_72_n_793

   PIN n_112099
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.634 0.0 59.662 0.163 ;
      END
   END n_112099

   PIN n_118917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.594 0.0 36.622 0.163 ;
      END
   END n_118917

   PIN n_119200
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.378 0.0 35.406 0.163 ;
      END
   END n_119200

   PIN n_122513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.93 0.0 66.958 0.163 ;
      END
   END n_122513

   PIN n_127504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.938 0.0 69.966 0.163 ;
      END
   END n_127504

   PIN n_127505
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.346 0.0 103.374 0.163 ;
      END
   END n_127505

   PIN n_137854
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.49 0.0 53.518 0.163 ;
      END
   END n_137854

   PIN n_140202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.226 0.0 130.254 0.163 ;
      END
   END n_140202

   PIN n_144103
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.25 0.0 43.278 0.163 ;
      END
   END n_144103

   PIN n_144157
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.058 0.0 43.086 0.163 ;
      END
   END n_144157

   PIN n_144176
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.794 0.0 23.822 0.163 ;
      END
   END n_144176

   PIN n_14438
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.49 0.0 29.518 0.163 ;
      END
   END n_14438

   PIN n_15497
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.658 0.0 4.686 0.163 ;
      END
   END n_15497

   PIN n_15502
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.362 0.0 29.39 0.163 ;
      END
   END n_15502

   PIN n_18035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.602 0.0 31.63 0.163 ;
      END
   END n_18035

   PIN n_19335
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.282 0.163 71.31 ;
      END
   END n_19335

   PIN n_19336
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.426 0.163 69.454 ;
      END
   END n_19336

   PIN n_19892
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.362 0.163 69.39 ;
      END
   END n_19892

   PIN n_20788
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.058 0.0 3.086 0.163 ;
      END
   END n_20788

   PIN n_20789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.994 0.0 3.022 0.163 ;
      END
   END n_20789

   PIN n_24618
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.322 0.163 78.35 ;
      END
   END n_24618

   PIN n_24620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.338 0.163 68.366 ;
      END
   END n_24620

   PIN n_24971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.498 0.0 128.526 0.163 ;
      END
   END n_24971

   PIN n_25653
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.09 0.0 135.118 0.163 ;
      END
   END n_25653

   PIN n_25723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.706 0.0 54.734 0.163 ;
      END
   END n_25723

   PIN n_25724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.026 0.0 55.054 0.163 ;
      END
   END n_25724

   PIN n_25959
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.066 0.0 70.094 0.163 ;
      END
   END n_25959

   PIN n_25961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.002 0.0 70.03 0.163 ;
      END
   END n_25961

   PIN n_26281
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.426 0.0 149.454 0.163 ;
      END
   END n_26281

   PIN n_26585
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.922 0.0 79.95 0.163 ;
      END
   END n_26585

   PIN n_26587
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.754 0.0 8.782 0.163 ;
      END
   END n_26587

   PIN n_26904
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.53 0.0 116.558 0.163 ;
      END
   END n_26904

   PIN n_26982
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 54.706 0.0 54.734 0.163 ;
      END
   END n_26982

   PIN n_27177
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.922 0.0 23.95 0.163 ;
      END
   END n_27177

   PIN n_27179
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.466 0.0 12.494 0.163 ;
      END
   END n_27179

   PIN n_27301
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.882 0.163 48.91 ;
      END
   END n_27301

   PIN n_27813
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.202 0.163 49.23 ;
      END
   END n_27813

   PIN n_27832
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.082 0.163 4.11 ;
      END
   END n_27832

   PIN n_27955
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.306 0.0 16.334 0.163 ;
      END
   END n_27955

   PIN n_27956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.242 0.0 16.27 0.163 ;
      END
   END n_27956

   PIN n_28339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.858 0.0 23.886 0.163 ;
      END
   END n_28339

   PIN n_28703
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.85 0.0 4.878 0.163 ;
      END
   END n_28703

   PIN n_29615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.13 0.163 102.158 ;
      END
   END n_29615

   PIN n_29657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.874 0.0 13.902 0.163 ;
      END
   END n_29657

   PIN n_29695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.074 0.0 73.102 0.163 ;
      END
   END n_29695

   PIN n_29942
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.714 0.0 73.742 0.163 ;
      END
   END n_29942

   PIN n_30391
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.434 0.0 16.462 0.163 ;
      END
   END n_30391

   PIN n_31042
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.106 0.0 5.134 0.163 ;
      END
   END n_31042

   PIN n_31230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.402 0.0 12.43 0.163 ;
      END
   END n_31230

   PIN n_34986
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.626 0.0 40.654 0.163 ;
      END
   END n_34986

   PIN n_35606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.018 0.0 20.046 0.163 ;
      END
   END n_35606

   PIN n_36793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.666 0.0 31.694 0.163 ;
      END
   END n_36793

   PIN n_37228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.674 0.0 50.702 0.163 ;
      END
   END n_37228

   PIN n_37268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.57 0.0 59.598 0.163 ;
      END
   END n_37268

   PIN n_37414
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.402 0.0 60.43 0.163 ;
      END
   END n_37414

   PIN n_37962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.442 0.0 35.47 0.163 ;
      END
   END n_37962

   PIN n_41276
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.026 0.163 7.054 ;
      END
   END n_41276

   PIN n_42685
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.626 0.0 40.654 0.163 ;
      END
   END n_42685

   PIN n_42686
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.562 0.0 40.59 0.163 ;
      END
   END n_42686

   PIN n_42769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.538 0.0 31.566 0.163 ;
      END
   END n_42769

   PIN n_43108
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.218 0.0 31.246 0.163 ;
      END
   END n_43108

   PIN n_49334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.426 0.163 45.454 ;
      END
   END n_49334

   PIN n_49644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.242 0.0 64.27 0.163 ;
      END
   END n_49644

   PIN n_52858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.186 0.0 43.214 0.163 ;
      END
   END n_52858

   PIN n_54999
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.314 0.0 35.342 0.163 ;
      END
   END n_54999

   PIN n_58856
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.026 0.0 39.054 0.163 ;
      END
   END n_58856

   PIN n_62942
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.442 0.0 75.47 0.163 ;
      END
   END n_62942

   PIN n_63427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.738 0.0 74.766 0.163 ;
      END
   END n_63427

   PIN n_65431
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.25 0.0 107.278 0.163 ;
      END
   END n_65431

   PIN n_65453
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.682 0.0 77.71 0.163 ;
      END
   END n_65453

   PIN n_65981
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.418 0.0 90.446 0.163 ;
      END
   END n_65981

   PIN n_66003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.042 0.0 93.07 0.163 ;
      END
   END n_66003

   PIN n_87308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.426 0.0 85.454 0.163 ;
      END
   END n_87308

   PIN n_87309
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.362 0.0 85.39 0.163 ;
      END
   END n_87309

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 158.72 106.24 ;
      LAYER V1 ;
         RECT 0.0 0.0 158.72 106.24 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 158.72 106.24 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 158.72 106.24 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 158.72 106.24 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 158.72 106.24 ;
      LAYER M1 ;
         RECT 0.0 0.0 158.72 106.24 ;
   END
END h4_mgc_matrix_mult_a

MACRO h3_mgc_matrix_mult_a
   CLASS BLOCK ;
   FOREIGN h3 ;
   ORIGIN 0 0 ;
   SIZE 154.688 BY 250.24 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN11777_n_66950
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.234 0.163 13.262 ;
      END
   END FE_OFN11777_n_66950

   PIN FE_OFN12461_n_66941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.562 0.082 40.59 ;
      END
   END FE_OFN12461_n_66941

   PIN FE_OFN12463_n_66941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.266 0.163 17.294 ;
      END
   END FE_OFN12463_n_66941

   PIN FE_OFN12466_n_66941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.666 0.163 55.694 ;
      END
   END FE_OFN12466_n_66941

   PIN FE_OFN12469_n_66941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.37 0.0 24.398 0.163 ;
      END
   END FE_OFN12469_n_66941

   PIN FE_OFN12475_n_66941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.762 0.0 35.79 0.163 ;
      END
   END FE_OFN12475_n_66941

   PIN FE_OFN12476_n_66941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.898 0.163 70.926 ;
      END
   END FE_OFN12476_n_66941

   PIN FE_OFN12505_n_66968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.578 0.163 78.606 ;
      END
   END FE_OFN12505_n_66968

   PIN FE_OFN12507_n_66968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.682 0.163 13.71 ;
      END
   END FE_OFN12507_n_66968

   PIN FE_OFN12512_n_66968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.954 0.0 19.982 0.163 ;
      END
   END FE_OFN12512_n_66968

   PIN FE_OFN12517_n_66968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.946 0.163 24.974 ;
      END
   END FE_OFN12517_n_66968

   PIN FE_OFN12520_n_66968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.722 0.163 36.75 ;
      END
   END FE_OFN12520_n_66968

   PIN FE_OFN12586_n_40826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.178 0.163 32.206 ;
      END
   END FE_OFN12586_n_40826

   PIN FE_OFN12925_n_66944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.402 0.0 20.43 0.163 ;
      END
   END FE_OFN12925_n_66944

   PIN FE_OFN12926_n_66944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.402 0.082 44.43 ;
      END
   END FE_OFN12926_n_66944

   PIN FE_OFN12929_n_66944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.17 0.082 21.198 ;
      END
   END FE_OFN12929_n_66944

   PIN FE_OFN13152_n_66961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.81 0.082 13.838 ;
      END
   END FE_OFN13152_n_66961

   PIN FE_OFN13959_n_40850
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.442 0.163 67.47 ;
      END
   END FE_OFN13959_n_40850

   PIN FE_OFN13962_n_40850
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.65 0.0 89.678 0.082 ;
      END
   END FE_OFN13962_n_40850

   PIN FE_OFN13963_n_40850
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.634 0.163 51.662 ;
      END
   END FE_OFN13963_n_40850

   PIN FE_OFN14315_n_67092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.266 0.0 129.294 0.163 ;
      END
   END FE_OFN14315_n_67092

   PIN FE_OFN14437_n_66941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.65 0.163 9.678 ;
      END
   END FE_OFN14437_n_66941

   PIN FE_OFN16001_n_66961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.97 0.163 1.998 ;
      END
   END FE_OFN16001_n_66961

   PIN FE_OFN17415_n_8277
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.346 0.163 63.374 ;
      END
   END FE_OFN17415_n_8277

   PIN FE_OFN4388_n_8279
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.842 0.163 97.87 ;
      END
   END FE_OFN4388_n_8279

   PIN FE_OFN4393_n_11208
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.874 0.163 93.902 ;
      END
   END FE_OFN4393_n_11208

   PIN FE_OFN4395_n_8397
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.098 0.163 90.126 ;
      END
   END FE_OFN4395_n_8397

   PIN FE_OFN4396_n_11207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 157.17 0.163 157.198 ;
      END
   END FE_OFN4396_n_11207

   PIN FE_OFN4457_n_9794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.258 0.163 86.286 ;
      END
   END FE_OFN4457_n_9794

   PIN FE_OFN4464_n_8278
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.522 0.163 105.55 ;
      END
   END FE_OFN4464_n_8278

   PIN FE_OFN4479_n_11214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.586 0.163 105.614 ;
      END
   END FE_OFN4479_n_11214

   PIN FE_OFN4483_n_11196
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 143.026 0.163 143.054 ;
      END
   END FE_OFN4483_n_11196

   PIN FE_OFN4485_n_8400
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 91.826 0.163 91.854 ;
      END
   END FE_OFN4485_n_8400

   PIN FE_OFN4487_n_8265
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.65 0.163 105.678 ;
      END
   END FE_OFN4487_n_8265

   PIN FE_OFN4489_n_8249
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.17 0.163 109.198 ;
      END
   END FE_OFN4489_n_8249

   PIN FE_OFN4531_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 134.642 0.163 134.67 ;
      END
   END FE_OFN4531_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_2_

   PIN FE_OFN4541_n_137715
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.49 0.163 117.518 ;
      END
   END FE_OFN4541_n_137715

   PIN FE_OFN5216_n_66958
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.842 0.163 57.87 ;
      END
   END FE_OFN5216_n_66958

   PIN FE_OFN5217_n_66958
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.874 0.163 5.902 ;
      END
   END FE_OFN5217_n_66958

   PIN FE_OFN5249_n_65559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 49.906 0.0 49.934 0.082 ;
      END
   END FE_OFN5249_n_65559

   PIN FE_OFN5641_delay_mul_ln34_unr6_unr7_stage2_stallmux_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 201.842 0.163 201.87 ;
      END
   END FE_OFN5641_delay_mul_ln34_unr6_unr7_stage2_stallmux_z_6_

   PIN FE_OFN8871_n_6526
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 220.658 0.163 220.686 ;
      END
   END FE_OFN8871_n_6526

   PIN FE_OFN8989_n_30545
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.946 250.077 8.974 250.24 ;
      END
   END FE_OFN8989_n_30545

   PIN FE_OFN9028_n_29931
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.09 250.077 31.118 250.24 ;
      END
   END FE_OFN9028_n_29931

   PIN FE_OFN9031_n_18065
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 232.306 0.163 232.334 ;
      END
   END FE_OFN9031_n_18065

   PIN FE_OFN9097_n_17577
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 213.042 0.163 213.07 ;
      END
   END FE_OFN9097_n_17577

   PIN delay_mul_ln34_unr4_unr8_stage2_stallmux_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 136.178 0.163 136.206 ;
      END
   END delay_mul_ln34_unr4_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr4_unr8_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.906 0.163 97.934 ;
      END
   END delay_mul_ln34_unr4_unr8_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr4_unr8_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.002 0.163 94.03 ;
      END
   END delay_mul_ln34_unr4_unr8_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr4_unr8_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.066 0.163 94.094 ;
      END
   END delay_mul_ln34_unr4_unr8_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr4_unr8_stage2_stallmux_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 120.882 0.163 120.91 ;
      END
   END delay_mul_ln34_unr4_unr8_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr4_unr8_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.234 0.163 109.262 ;
      END
   END delay_mul_ln34_unr4_unr8_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr4_unr8_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.554 0.163 101.582 ;
      END
   END delay_mul_ln34_unr4_unr8_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 132.402 0.163 132.43 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr5_unr4_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 147.762 0.163 147.79 ;
      END
   END delay_mul_ln34_unr5_unr4_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr5_unr4_stage2_stallmux_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 155.314 0.163 155.342 ;
      END
   END delay_mul_ln34_unr5_unr4_stage2_stallmux_z_14_

   PIN n_100713
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.41 0.163 55.438 ;
      END
   END n_100713

   PIN n_100723
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.146 0.163 44.174 ;
      END
   END n_100723

   PIN n_100936
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 124.722 0.163 124.75 ;
      END
   END n_100936

   PIN n_103466
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.93 0.163 66.958 ;
      END
   END n_103466

   PIN n_103926
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.706 0.163 102.734 ;
      END
   END n_103926

   PIN n_104085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 124.786 0.163 124.814 ;
      END
   END n_104085

   PIN n_104088
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 128.498 0.163 128.526 ;
      END
   END n_104088

   PIN n_106337
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.578 0.0 62.606 0.163 ;
      END
   END n_106337

   PIN n_107599
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 129.01 0.163 129.038 ;
      END
   END n_107599

   PIN n_108566
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.618 0.163 101.646 ;
      END
   END n_108566

   PIN n_108600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 132.466 0.163 132.494 ;
      END
   END n_108600

   PIN n_109675
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.818 0.0 56.846 0.163 ;
      END
   END n_109675

   PIN n_110044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.61 0.163 82.638 ;
      END
   END n_110044

   PIN n_110200
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.298 0.163 109.326 ;
      END
   END n_110200

   PIN n_111224
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 84.722 0.163 84.75 ;
      END
   END n_111224

   PIN n_111289
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.482 0.163 82.51 ;
      END
   END n_111289

   PIN n_137850
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 139.762 0.163 139.79 ;
      END
   END n_137850

   PIN n_14225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 128.434 0.163 128.462 ;
      END
   END n_14225

   PIN n_14437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.314 250.077 11.342 250.24 ;
      END
   END n_14437

   PIN n_17579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 224.626 0.163 224.654 ;
      END
   END n_17579

   PIN n_17740
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.554 0.163 117.582 ;
      END
   END n_17740

   PIN n_19137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 129.586 0.163 129.614 ;
      END
   END n_19137

   PIN n_19430
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.362 0.163 109.39 ;
      END
   END n_19430

   PIN n_21697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 220.722 0.163 220.75 ;
      END
   END n_21697

   PIN n_22575
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 192.242 0.163 192.27 ;
      END
   END n_22575

   PIN n_22812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 237.042 0.163 237.07 ;
      END
   END n_22812

   PIN n_22823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 247.602 0.163 247.63 ;
      END
   END n_22823

   PIN n_23106
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.322 0.163 86.35 ;
      END
   END n_23106

   PIN n_23397
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 218.546 0.163 218.574 ;
      END
   END n_23397

   PIN n_24070
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 213.106 0.163 213.134 ;
      END
   END n_24070

   PIN n_24076
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.026 250.077 55.054 250.24 ;
      END
   END n_24076

   PIN n_24694
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 213.17 0.163 213.198 ;
      END
   END n_24694

   PIN n_25002
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 209.202 0.163 209.23 ;
      END
   END n_25002

   PIN n_25685
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 205.426 0.163 205.454 ;
      END
   END n_25685

   PIN n_25764
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 164.786 0.163 164.814 ;
      END
   END n_25764

   PIN n_26319
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 173.746 0.163 173.774 ;
      END
   END n_26319

   PIN n_27216
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 224.562 0.163 224.59 ;
      END
   END n_27216

   PIN n_30014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 236.402 0.163 236.43 ;
      END
   END n_30014

   PIN n_4303
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.81 0.163 93.838 ;
      END
   END n_4303

   PIN n_66951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.682 0.163 5.71 ;
      END
   END n_66951

   PIN n_67661
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.794 0.163 47.822 ;
      END
   END n_67661

   PIN n_68032
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.794 0.163 31.822 ;
      END
   END n_68032

   PIN n_68033
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.73 0.163 31.758 ;
      END
   END n_68033

   PIN n_69311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.498 0.0 24.526 0.163 ;
      END
   END n_69311

   PIN n_72597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.178 0.0 24.206 0.163 ;
      END
   END n_72597

   PIN n_72604
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.962 0.163 30.99 ;
      END
   END n_72604

   PIN n_72605
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.218 0.163 31.246 ;
      END
   END n_72605

   PIN n_72988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.178 0.163 40.206 ;
      END
   END n_72988

   PIN n_72992
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.594 0.163 28.622 ;
      END
   END n_72992

   PIN n_72993
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.658 0.163 28.686 ;
      END
   END n_72993

   PIN n_73152
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.146 0.0 28.174 0.163 ;
      END
   END n_73152

   PIN n_73468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.866 0.0 58.894 0.163 ;
      END
   END n_73468

   PIN n_73744
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.538 0.163 55.566 ;
      END
   END n_73744

   PIN n_73917
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.434 0.0 24.462 0.163 ;
      END
   END n_73917

   PIN n_73948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.986 0.163 24.014 ;
      END
   END n_73948

   PIN n_74101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.282 0.163 63.31 ;
      END
   END n_74101

   PIN n_74594
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.242 0.0 24.27 0.163 ;
      END
   END n_74594

   PIN n_75501
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.05 0.163 24.078 ;
      END
   END n_75501

   PIN n_75780
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.89 0.0 11.918 0.163 ;
      END
   END n_75780

   PIN n_75876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.762 0.163 75.79 ;
      END
   END n_75876

   PIN n_76534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.93 0.0 50.958 0.163 ;
      END
   END n_76534

   PIN n_79296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.178 0.0 40.206 0.163 ;
      END
   END n_79296

   PIN n_79300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.618 0.0 45.646 0.163 ;
      END
   END n_79300

   PIN n_79437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.922 0.163 23.95 ;
      END
   END n_79437

   PIN n_79786
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.194 0.0 62.222 0.163 ;
      END
   END n_79786

   PIN n_79790
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.146 0.163 36.174 ;
      END
   END n_79790

   PIN n_80033
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.498 0.0 152.526 0.163 ;
      END
   END n_80033

   PIN n_80045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.026 0.0 39.054 0.163 ;
      END
   END n_80045

   PIN n_80047
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.898 0.0 54.926 0.163 ;
      END
   END n_80047

   PIN n_80051
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.306 0.0 120.334 0.163 ;
      END
   END n_80051

   PIN n_81552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.242 0.163 48.27 ;
      END
   END n_81552

   PIN n_81553
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.962 0.163 46.99 ;
      END
   END n_81553

   PIN n_81623
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.258 0.0 62.286 0.163 ;
      END
   END n_81623

   PIN n_81655
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.714 0.0 33.742 0.163 ;
      END
   END n_81655

   PIN n_81678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.802 0.0 58.83 0.163 ;
      END
   END n_81678

   PIN n_81735
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.242 0.0 120.27 0.163 ;
      END
   END n_81735

   PIN n_82059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.082 0.163 36.11 ;
      END
   END n_82059

   PIN n_82060
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.21 0.163 36.238 ;
      END
   END n_82060

   PIN n_82522
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.162 0.163 90.19 ;
      END
   END n_82522

   PIN n_82528
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.546 0.163 82.574 ;
      END
   END n_82528

   PIN n_82532
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.082 0.163 4.11 ;
      END
   END n_82532

   PIN n_82968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.858 0.163 47.886 ;
      END
   END n_82968

   PIN n_86363
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.042 0.0 29.07 0.163 ;
      END
   END n_86363

   PIN n_86802
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.57 0.0 83.598 0.163 ;
      END
   END n_86802

   PIN n_87172
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.962 0.0 54.99 0.163 ;
      END
   END n_87172

   PIN n_87450
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.586 0.0 57.614 0.163 ;
      END
   END n_87450

   PIN n_87451
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.522 0.0 49.55 0.163 ;
      END
   END n_87451

   PIN n_87971
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.698 0.163 51.726 ;
      END
   END n_87971

   PIN n_88095
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.042 0.163 77.07 ;
      END
   END n_88095

   PIN n_88096
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.106 0.163 77.134 ;
      END
   END n_88096

   PIN n_88390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.586 0.163 9.614 ;
      END
   END n_88390

   PIN n_89684
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.818 0.0 96.846 0.163 ;
      END
   END n_89684

   PIN n_89697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.194 0.0 78.222 0.163 ;
      END
   END n_89697

   PIN n_89726
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.546 0.0 42.574 0.163 ;
      END
   END n_89726

   PIN n_89763
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.546 0.0 114.574 0.163 ;
      END
   END n_89763

   PIN n_90132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.474 0.163 55.502 ;
      END
   END n_90132

   PIN n_90144
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.666 0.163 47.694 ;
      END
   END n_90144

   PIN n_90579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.938 0.163 93.966 ;
      END
   END n_90579

   PIN n_91470
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.45 0.0 62.478 0.163 ;
      END
   END n_91470

   PIN n_91617
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.674 0.0 50.702 0.163 ;
      END
   END n_91617

   PIN n_92981
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.458 0.0 89.486 0.163 ;
      END
   END n_92981

   PIN n_93705
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.162 0.0 74.19 0.163 ;
      END
   END n_93705

   PIN n_94165
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.506 0.0 75.534 0.163 ;
      END
   END n_94165

   PIN n_94212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.122 0.0 107.15 0.163 ;
      END
   END n_94212

   PIN n_94213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.37 0.0 112.398 0.163 ;
      END
   END n_94213

   PIN n_94385
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.57 0.163 51.598 ;
      END
   END n_94385

   PIN n_94604
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.386 0.163 94.414 ;
      END
   END n_94604

   PIN n_95206
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.482 0.0 42.51 0.163 ;
      END
   END n_95206

   PIN n_96024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.762 0.0 131.79 0.163 ;
      END
   END n_96024

   PIN n_96027
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.018 0.0 132.046 0.163 ;
      END
   END n_96027

   PIN n_96606
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.226 0.163 90.254 ;
      END
   END n_96606

   PIN n_99922
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.802 0.163 66.83 ;
      END
   END n_99922

   PIN FE_OFN11773_n_66950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.642 0.163 22.67 ;
      END
   END FE_OFN11773_n_66950

   PIN FE_OFN11776_n_66950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.474 0.0 39.502 0.082 ;
      END
   END FE_OFN11776_n_66950

   PIN FE_OFN11782_n_66950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.738 0.0 58.766 0.163 ;
      END
   END FE_OFN11782_n_66950

   PIN FE_OFN11785_n_66950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.306 0.0 24.334 0.082 ;
      END
   END FE_OFN11785_n_66950

   PIN FE_OFN12151_n_40871
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.674 0.0 58.702 0.082 ;
      END
   END FE_OFN12151_n_40871

   PIN FE_OFN12262_n_66958
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.042 0.163 21.07 ;
      END
   END FE_OFN12262_n_66958

   PIN FE_OFN12456_n_66941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.658 0.163 36.686 ;
      END
   END FE_OFN12456_n_66941

   PIN FE_OFN12462_n_66941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.81 0.163 5.838 ;
      END
   END FE_OFN12462_n_66941

   PIN FE_OFN12464_n_66941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.402 0.163 36.43 ;
      END
   END FE_OFN12464_n_66941

   PIN FE_OFN12470_n_66941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 36.466 0.163 36.494 ;
      END
   END FE_OFN12470_n_66941

   PIN FE_OFN12500_n_66968
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.978 0.163 29.006 ;
      END
   END FE_OFN12500_n_66968

   PIN FE_OFN12502_n_66968
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.322 0.163 14.35 ;
      END
   END FE_OFN12502_n_66968

   PIN FE_OFN12514_n_66968
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.202 0.163 17.23 ;
      END
   END FE_OFN12514_n_66968

   PIN FE_OFN12581_n_40826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.658 0.0 36.686 0.163 ;
      END
   END FE_OFN12581_n_40826

   PIN FE_OFN12591_n_40826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.602 0.0 39.63 0.082 ;
      END
   END FE_OFN12591_n_40826

   PIN FE_OFN12593_n_40826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.978 0.163 21.006 ;
      END
   END FE_OFN12593_n_40826

   PIN FE_OFN12915_n_66944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.906 0.163 1.934 ;
      END
   END FE_OFN12915_n_66944

   PIN FE_OFN12919_n_66944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.322 0.163 22.35 ;
      END
   END FE_OFN12919_n_66944

   PIN FE_OFN12943_n_67234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 32.37 0.082 32.398 ;
      END
   END FE_OFN12943_n_67234

   PIN FE_OFN13149_n_66961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.85 0.163 20.878 ;
      END
   END FE_OFN13149_n_66961

   PIN FE_OFN13155_n_66961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.93 0.0 58.958 0.082 ;
      END
   END FE_OFN13155_n_66961

   PIN FE_OFN13156_n_66961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.082 0.082 68.11 ;
      END
   END FE_OFN13156_n_66961

   PIN FE_OFN13160_n_66961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.786 0.163 20.814 ;
      END
   END FE_OFN13160_n_66961

   PIN FE_OFN13177_n_67154
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.034 0.163 2.062 ;
      END
   END FE_OFN13177_n_67154

   PIN FE_OFN13643_n_40808
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.042 0.163 13.07 ;
      END
   END FE_OFN13643_n_40808

   PIN FE_OFN13953_n_40848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.338 0.163 36.366 ;
      END
   END FE_OFN13953_n_40848

   PIN FE_OFN13957_n_40849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.202 0.163 57.23 ;
      END
   END FE_OFN13957_n_40849

   PIN FE_OFN13969_n_40851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.026 0.082 71.054 ;
      END
   END FE_OFN13969_n_40851

   PIN FE_OFN14037_n_40809
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 76.082 0.163 76.11 ;
      END
   END FE_OFN14037_n_40809

   PIN FE_OFN14042_n_40810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.802 0.163 74.83 ;
      END
   END FE_OFN14042_n_40810

   PIN FE_OFN14064_n_67235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.546 0.163 18.574 ;
      END
   END FE_OFN14064_n_67235

   PIN FE_OFN14067_n_67237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.882 0.163 24.91 ;
      END
   END FE_OFN14067_n_67237

   PIN FE_OFN14094_n_67196
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.33 0.163 17.358 ;
      END
   END FE_OFN14094_n_67196

   PIN FE_OFN14100_n_40807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.282 0.0 47.31 0.163 ;
      END
   END FE_OFN14100_n_40807

   PIN FE_OFN14313_n_67092
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.33 0.0 129.358 0.163 ;
      END
   END FE_OFN14313_n_67092

   PIN FE_OFN14354_n_65559
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.274 0.163 36.302 ;
      END
   END FE_OFN14354_n_65559

   PIN FE_OFN14377_n_67149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 21.106 0.163 21.134 ;
      END
   END FE_OFN14377_n_67149

   PIN FE_OFN14439_n_66941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.274 0.163 44.302 ;
      END
   END FE_OFN14439_n_66941

   PIN FE_OFN14502_n_40871
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.05 0.082 40.078 ;
      END
   END FE_OFN14502_n_40871

   PIN FE_OFN15991_n_65559
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.946 0.163 40.974 ;
      END
   END FE_OFN15991_n_65559

   PIN FE_OFN15996_n_66956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.042 0.163 29.07 ;
      END
   END FE_OFN15996_n_66956

   PIN FE_OFN17405_n_9785
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 218.482 0.163 218.51 ;
      END
   END FE_OFN17405_n_9785

   PIN FE_OFN17406_n_11207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 166.002 0.163 166.03 ;
      END
   END FE_OFN17406_n_11207

   PIN FE_OFN17421_n_8265
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 142.962 0.163 142.99 ;
      END
   END FE_OFN17421_n_8265

   PIN FE_OFN17424_delay_mul_ln34_unr4_unr8_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 182.258 0.163 182.286 ;
      END
   END FE_OFN17424_delay_mul_ln34_unr4_unr8_stage2_stallmux_z_4_

   PIN FE_OFN17454_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 150.642 0.163 150.67 ;
      END
   END FE_OFN17454_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_2_

   PIN FE_OFN19163_n_8279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 193.522 0.163 193.55 ;
      END
   END FE_OFN19163_n_8279

   PIN FE_OFN4392_n_11208
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 120.562 0.163 120.59 ;
      END
   END FE_OFN4392_n_11208

   PIN FE_OFN4394_n_8397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 100.146 0.163 100.174 ;
      END
   END FE_OFN4394_n_8397

   PIN FE_OFN4478_n_11214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.106 0.163 109.134 ;
      END
   END FE_OFN4478_n_11214

   PIN FE_OFN4484_n_8400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 91.762 0.163 91.79 ;
      END
   END FE_OFN4484_n_8400

   PIN FE_OFN4488_n_8249
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.042 0.163 109.07 ;
      END
   END FE_OFN4488_n_8249

   PIN FE_OFN4522_delay_mul_ln34_unr4_unr8_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 173.682 0.163 173.71 ;
      END
   END FE_OFN4522_delay_mul_ln34_unr4_unr8_stage2_stallmux_z_2_

   PIN FE_OFN4540_n_137715
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.426 0.163 117.454 ;
      END
   END FE_OFN4540_n_137715

   PIN FE_OFN5096_n_66960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.874 0.0 77.902 0.082 ;
      END
   END FE_OFN5096_n_66960

   PIN FE_OFN5273_n_40871
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.346 0.0 47.374 0.082 ;
      END
   END FE_OFN5273_n_40871

   PIN FE_OFN5289_n_66950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.09 0.082 31.118 ;
      END
   END FE_OFN5289_n_66950

   PIN FE_OFN5335_n_66955
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.082 0.163 44.11 ;
      END
   END FE_OFN5335_n_66955

   PIN FE_OFN5339_n_66955
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.922 0.163 39.95 ;
      END
   END FE_OFN5339_n_66955

   PIN FE_OFN5388_n_66961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.722 0.0 12.75 0.163 ;
      END
   END FE_OFN5388_n_66961

   PIN FE_OFN5455_n_67234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.842 0.163 1.87 ;
      END
   END FE_OFN5455_n_67234

   PIN FE_OFN5517_n_67154
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.914 0.163 20.942 ;
      END
   END FE_OFN5517_n_67154

   PIN FE_OFN5522_n_67150
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.818 0.163 24.846 ;
      END
   END FE_OFN5522_n_67150

   PIN FE_OFN5557_n_67036
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.218 0.0 47.246 0.163 ;
      END
   END FE_OFN5557_n_67036

   PIN FE_OFN9027_n_29931
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 174.642 0.163 174.67 ;
      END
   END FE_OFN9027_n_29931

   PIN FE_OFN9806_b_5_5_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.306 0.163 32.334 ;
      END
   END FE_OFN9806_b_5_5_1

   PIN b_5_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.602 0.082 31.63 ;
      END
   END b_5_3_0

   PIN b_5_3_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.882 0.082 48.91 ;
      END
   END b_5_3_1

   PIN b_5_3_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.162 0.082 50.19 ;
      END
   END b_5_3_5

   PIN b_5_3_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.73 0.163 47.758 ;
      END
   END b_5_3_6

   PIN b_5_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.606 67.122 154.688 67.15 ;
      END
   END b_5_4_0

   PIN b_5_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.606 47.922 154.688 47.95 ;
      END
   END b_5_4_1

   PIN b_5_4_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.525 82.546 154.688 82.574 ;
      END
   END b_5_4_10

   PIN b_5_4_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.525 71.09 154.688 71.118 ;
      END
   END b_5_4_11

   PIN b_5_4_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.525 78.77 154.688 78.798 ;
      END
   END b_5_4_12

   PIN b_5_4_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.525 71.026 154.688 71.054 ;
      END
   END b_5_4_13

   PIN b_5_4_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.525 70.962 154.688 70.99 ;
      END
   END b_5_4_14

   PIN b_5_4_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.45 0.082 22.478 ;
      END
   END b_5_4_2

   PIN b_5_4_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.57 0.082 67.598 ;
      END
   END b_5_4_3

   PIN b_5_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.514 0.0 78.542 0.082 ;
      END
   END b_5_4_4

   PIN b_5_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.606 74.802 154.688 74.83 ;
      END
   END b_5_4_5

   PIN b_5_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.525 94.066 154.688 94.094 ;
      END
   END b_5_4_6

   PIN b_5_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.106 0.163 13.134 ;
      END
   END b_5_4_7

   PIN b_5_4_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.194 0.0 46.222 0.163 ;
      END
   END b_5_4_8

   PIN b_5_4_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.525 86.386 154.688 86.414 ;
      END
   END b_5_4_9

   PIN b_5_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 142.194 0.0 142.222 0.082 ;
      END
   END b_5_6_0

   PIN b_5_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.946 0.0 120.974 0.082 ;
      END
   END b_5_6_1

   PIN b_5_6_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.525 55.666 154.688 55.694 ;
      END
   END b_5_6_10

   PIN b_5_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.606 28.722 154.688 28.75 ;
      END
   END b_5_6_2

   PIN b_5_6_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.018 0.0 52.046 0.082 ;
      END
   END b_5_6_3

   PIN b_5_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.186 0.0 51.214 0.082 ;
      END
   END b_5_6_4

   PIN b_5_6_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 154.606 82.162 154.688 82.19 ;
      END
   END b_5_6_5

   PIN b_5_6_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.626 0.0 48.654 0.163 ;
      END
   END b_5_6_6

   PIN b_5_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.482 0.0 82.51 0.163 ;
      END
   END b_5_6_7

   PIN b_5_6_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.746 0.0 45.774 0.163 ;
      END
   END b_5_6_8

   PIN b_5_6_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.33 0.0 65.358 0.163 ;
      END
   END b_5_6_9

   PIN b_5_9_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.346 0.082 31.374 ;
      END
   END b_5_9_0

   PIN b_5_9_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.602 0.163 47.63 ;
      END
   END b_5_9_1

   PIN b_5_9_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.786 0.082 28.814 ;
      END
   END b_5_9_2

   PIN delay_mul_ln34_unr3_unr8_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.13 0.0 38.158 0.163 ;
      END
   END delay_mul_ln34_unr3_unr8_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 196.082 0.163 196.11 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 246.002 0.163 246.03 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 212.978 0.163 213.006 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_q_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 218.482 0.163 218.51 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_q_3_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 190.002 0.163 190.03 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 157.106 0.163 157.134 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr4_unr8_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 146.802 0.163 146.83 ;
      END
   END delay_mul_ln34_unr4_unr8_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr5_unr5_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.594 0.163 36.622 ;
      END
   END delay_mul_ln34_unr5_unr5_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr5_unr5_stage2_stallmux_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.522 0.163 65.55 ;
      END
   END delay_mul_ln34_unr5_unr5_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr5_unr5_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.994 0.163 67.022 ;
      END
   END delay_mul_ln34_unr5_unr5_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr5_unr5_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.242 0.163 32.27 ;
      END
   END delay_mul_ln34_unr5_unr5_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr5_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.434 0.163 40.462 ;
      END
   END delay_mul_ln34_unr5_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr5_unr8_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.746 0.163 5.774 ;
      END
   END delay_mul_ln34_unr5_unr8_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr5_unr8_stage2_stallmux_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 125.682 0.163 125.71 ;
      END
   END delay_mul_ln34_unr5_unr8_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr6_unr3_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 219.186 0.163 219.214 ;
      END
   END delay_mul_ln34_unr6_unr3_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr6_unr7_stage2_stallmux_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 205.362 0.163 205.39 ;
      END
   END delay_mul_ln34_unr6_unr7_stage2_stallmux_z_6_

   PIN delay_mul_ln34_unr6_unr8_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 179.442 0.163 179.47 ;
      END
   END delay_mul_ln34_unr6_unr8_stage2_stallmux_q_15_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 183.602 0.082 183.63 ;
      END
   END ispd_clk

   PIN n_100719
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.826 0.163 51.854 ;
      END
   END n_100719

   PIN n_100722
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.018 0.163 44.046 ;
      END
   END n_100722

   PIN n_101748
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.866 0.163 66.894 ;
      END
   END n_101748

   PIN n_103932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.21 0.163 44.238 ;
      END
   END n_103932

   PIN n_104087
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 128.946 0.163 128.974 ;
      END
   END n_104087

   PIN n_10440
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 156.402 0.163 156.43 ;
      END
   END n_10440

   PIN n_105093
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.026 0.0 55.054 0.163 ;
      END
   END n_105093

   PIN n_105235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.73 0.163 55.758 ;
      END
   END n_105235

   PIN n_105237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.218 0.163 71.246 ;
      END
   END n_105237

   PIN n_106469
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.41 0.163 63.438 ;
      END
   END n_106469

   PIN n_106554
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 128.882 0.163 128.91 ;
      END
   END n_106554

   PIN n_108572
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 51.826 0.163 51.854 ;
      END
   END n_108572

   PIN n_110944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 111.602 0.163 111.63 ;
      END
   END n_110944

   PIN n_110947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 132.53 0.163 132.558 ;
      END
   END n_110947

   PIN n_11196
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 164.722 0.163 164.75 ;
      END
   END n_11196

   PIN n_12058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 137.906 0.163 137.934 ;
      END
   END n_12058

   PIN n_12059
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 137.842 0.163 137.87 ;
      END
   END n_12059

   PIN n_13500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.97 0.0 17.998 0.163 ;
      END
   END n_13500

   PIN n_137713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 228.402 0.163 228.43 ;
      END
   END n_137713

   PIN n_137779
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 209.522 0.163 209.55 ;
      END
   END n_137779

   PIN n_137786
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 147.442 0.163 147.47 ;
      END
   END n_137786

   PIN n_137843
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 228.082 0.163 228.11 ;
      END
   END n_137843

   PIN n_137880
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 236.018 0.163 236.046 ;
      END
   END n_137880

   PIN n_143962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.37 0.163 40.398 ;
      END
   END n_143962

   PIN n_144202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.21 0.0 36.238 0.163 ;
      END
   END n_144202

   PIN n_16583
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 120.946 0.163 120.974 ;
      END
   END n_16583

   PIN n_17577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 210.802 0.163 210.83 ;
      END
   END n_17577

   PIN n_17741
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.362 0.163 117.39 ;
      END
   END n_17741

   PIN n_18065
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 186.226 0.163 186.254 ;
      END
   END n_18065

   PIN n_18390
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 186.162 0.163 186.19 ;
      END
   END n_18390

   PIN n_19302
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.786 0.0 12.814 0.163 ;
      END
   END n_19302

   PIN n_20628
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.882 0.0 16.91 0.163 ;
      END
   END n_20628

   PIN n_21700
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.994 0.0 27.022 0.163 ;
      END
   END n_21700

   PIN n_22237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 157.042 0.163 157.07 ;
      END
   END n_22237

   PIN n_22437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 182.962 0.163 182.99 ;
      END
   END n_22437

   PIN n_22574
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 186.29 0.163 186.318 ;
      END
   END n_22574

   PIN n_22713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 156.722 0.163 156.75 ;
      END
   END n_22713

   PIN n_23320
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 191.602 0.163 191.63 ;
      END
   END n_23320

   PIN n_23322
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 193.842 0.163 193.87 ;
      END
   END n_23322

   PIN n_23688
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.386 0.163 86.414 ;
      END
   END n_23688

   PIN n_24904
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.13 0.163 94.158 ;
      END
   END n_24904

   PIN n_24905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.154 0.163 71.182 ;
      END
   END n_24905

   PIN n_25939
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 165.362 0.163 165.39 ;
      END
   END n_25939

   PIN n_26597
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 201.202 0.163 201.23 ;
      END
   END n_26597

   PIN n_29601
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 236.722 0.163 236.75 ;
      END
   END n_29601

   PIN n_30545
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.314 250.077 3.342 250.24 ;
      END
   END n_30545

   PIN n_41482
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.218 0.0 47.246 0.163 ;
      END
   END n_41482

   PIN n_41492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.418 0.0 66.446 0.163 ;
      END
   END n_41492

   PIN n_41540
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.218 0.163 63.246 ;
      END
   END n_41540

   PIN n_4506
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 129.522 0.163 129.55 ;
      END
   END n_4506

   PIN n_4623
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 219.122 0.163 219.15 ;
      END
   END n_4623

   PIN n_6549
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 227.442 0.163 227.47 ;
      END
   END n_6549

   PIN n_66953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.882 0.163 32.91 ;
      END
   END n_66953

   PIN n_66956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 32.114 0.082 32.142 ;
      END
   END n_66956

   PIN n_66959
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.482 0.082 58.51 ;
      END
   END n_66959

   PIN n_67155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.89 0.163 43.918 ;
      END
   END n_67155

   PIN n_67235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.986 0.163 32.014 ;
      END
   END n_67235

   PIN n_67643
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.53 0.163 36.558 ;
      END
   END n_67643

   PIN n_68016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.562 0.163 56.59 ;
      END
   END n_68016

   PIN n_70069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.522 0.163 9.55 ;
      END
   END n_70069

   PIN n_72452
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.826 0.163 43.854 ;
      END
   END n_72452

   PIN n_72987
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.642 0.163 38.67 ;
      END
   END n_72987

   PIN n_73547
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.906 0.163 57.934 ;
      END
   END n_73547

   PIN n_73658
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.034 0.163 90.062 ;
      END
   END n_73658

   PIN n_73743
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.602 0.163 55.63 ;
      END
   END n_73743

   PIN n_75140
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.698 0.0 35.726 0.163 ;
      END
   END n_75140

   PIN n_75485
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.386 0.0 70.414 0.163 ;
      END
   END n_75485

   PIN n_75486
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.274 0.0 68.302 0.163 ;
      END
   END n_75486

   PIN n_76729
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.146 0.0 124.174 0.163 ;
      END
   END n_76729

   PIN n_76730
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.386 0.0 118.414 0.163 ;
      END
   END n_76730

   PIN n_77155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.306 0.0 24.334 0.163 ;
      END
   END n_77155

   PIN n_77156
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.994 0.0 59.022 0.163 ;
      END
   END n_77156

   PIN n_77250
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.394 0.0 113.422 0.163 ;
      END
   END n_77250

   PIN n_81656
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.522 0.0 33.55 0.163 ;
      END
   END n_81656

   PIN n_82074
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.914 0.163 28.942 ;
      END
   END n_82074

   PIN n_8277
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 100.082 0.163 100.11 ;
      END
   END n_8277

   PIN n_8278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 170.866 0.163 170.894 ;
      END
   END n_8278

   PIN n_83010
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.466 0.163 36.494 ;
      END
   END n_83010

   PIN n_86823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.482 0.163 66.51 ;
      END
   END n_86823

   PIN n_86974
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.89 0.163 51.918 ;
      END
   END n_86974

   PIN n_89835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.922 0.0 127.95 0.163 ;
      END
   END n_89835

   PIN n_90145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.842 0.163 41.87 ;
      END
   END n_90145

   PIN n_90146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.954 0.163 43.982 ;
      END
   END n_90146

   PIN n_90147
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.074 0.163 49.102 ;
      END
   END n_90147

   PIN n_90149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.33 0.163 49.358 ;
      END
   END n_90149

   PIN n_90158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.53 0.163 44.558 ;
      END
   END n_90158

   PIN n_91623
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.322 0.163 94.35 ;
      END
   END n_91623

   PIN n_93661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.786 0.163 36.814 ;
      END
   END n_93661

   PIN n_94379
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.01 0.163 49.038 ;
      END
   END n_94379

   PIN n_95186
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.306 0.163 40.334 ;
      END
   END n_95186

   PIN n_95187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.242 0.163 40.27 ;
      END
   END n_95187

   PIN n_96274
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 45.426 0.163 45.454 ;
      END
   END n_96274

   PIN n_9777
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 140.082 0.163 140.11 ;
      END
   END n_9777

   PIN n_9778
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 138.482 0.163 138.51 ;
      END
   END n_9778

   PIN n_9794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.642 0.163 102.67 ;
      END
   END n_9794

   PIN n_98566
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.762 0.163 51.79 ;
      END
   END n_98566

   PIN n_98772
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.642 0.163 78.67 ;
      END
   END n_98772

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 154.688 250.24 ;
      LAYER V1 ;
         RECT 0.0 0.0 154.688 250.24 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 154.688 250.24 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 154.688 250.24 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 154.688 250.24 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 154.688 250.24 ;
      LAYER M1 ;
         RECT 0.0 0.0 154.688 250.24 ;
   END
END h3_mgc_matrix_mult_a

MACRO h2_mgc_matrix_mult_a
   CLASS BLOCK ;
   FOREIGN h2 ;
   ORIGIN 0 0 ;
   SIZE 249.792 BY 117.76 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN10016_b_4_4_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.154 0.0 55.182 0.163 ;
      END
   END FE_OFN10016_b_4_4_7

   PIN FE_OFN10107_b_4_2_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.338 0.0 60.366 0.163 ;
      END
   END FE_OFN10107_b_4_2_1

   PIN FE_OFN11689_n_140213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 76.914 249.792 76.942 ;
      END
   END FE_OFN11689_n_140213

   PIN FE_OFN11938_n_142850
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.986 0.0 96.014 0.163 ;
      END
   END FE_OFN11938_n_142850

   PIN FE_OFN12338_n_41013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.522 249.792 41.55 ;
      END
   END FE_OFN12338_n_41013

   PIN FE_OFN12341_n_41013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.746 249.792 29.774 ;
      END
   END FE_OFN12341_n_41013

   PIN FE_OFN12622_n_143670
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 36.978 249.792 37.006 ;
      END
   END FE_OFN12622_n_143670

   PIN FE_OFN12767_n_41734
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.498 249.792 40.526 ;
      END
   END FE_OFN12767_n_41734

   PIN FE_OFN12972_n_41962
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 225.394 0.0 225.422 0.163 ;
      END
   END FE_OFN12972_n_41962

   PIN FE_OFN13039_n_40828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.386 249.792 14.414 ;
      END
   END FE_OFN13039_n_40828

   PIN FE_OFN13195_n_137475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.45 249.792 14.478 ;
      END
   END FE_OFN13195_n_137475

   PIN FE_OFN13196_n_137475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.562 249.792 32.59 ;
      END
   END FE_OFN13196_n_137475

   PIN FE_OFN13200_n_137235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.314 249.792 11.342 ;
      END
   END FE_OFN13200_n_137235

   PIN FE_OFN13211_n_143630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 25.266 249.792 25.294 ;
      END
   END FE_OFN13211_n_143630

   PIN FE_OFN13228_n_143481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 189.106 0.0 189.134 0.163 ;
      END
   END FE_OFN13228_n_143481

   PIN FE_OFN13229_n_143481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 44.786 249.792 44.814 ;
      END
   END FE_OFN13229_n_143481

   PIN FE_OFN13244_n_41374
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 203.634 0.0 203.662 0.163 ;
      END
   END FE_OFN13244_n_41374

   PIN FE_OFN13247_n_143370
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.202 249.792 33.23 ;
      END
   END FE_OFN13247_n_143370

   PIN FE_OFN13354_n_41014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.602 249.792 55.63 ;
      END
   END FE_OFN13354_n_41014

   PIN FE_OFN13387_n_41612
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 28.85 249.792 28.878 ;
      END
   END FE_OFN13387_n_41612

   PIN FE_OFN13390_n_41612
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.626 249.792 32.654 ;
      END
   END FE_OFN13390_n_41612

   PIN FE_OFN13420_n_41709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.554 249.792 21.582 ;
      END
   END FE_OFN13420_n_41709

   PIN FE_OFN13421_n_41709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 10.866 249.792 10.894 ;
      END
   END FE_OFN13421_n_41709

   PIN FE_OFN13527_n_137233
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 13.938 249.792 13.966 ;
      END
   END FE_OFN13527_n_137233

   PIN FE_OFN13530_n_137233
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.162 0.0 242.19 0.163 ;
      END
   END FE_OFN13530_n_137233

   PIN FE_OFN13619_n_41963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.618 249.792 21.646 ;
      END
   END FE_OFN13619_n_41963

   PIN FE_OFN13620_n_41963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 202.226 0.0 202.254 0.163 ;
      END
   END FE_OFN13620_n_41963

   PIN FE_OFN13621_n_41963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.426 249.792 37.454 ;
      END
   END FE_OFN13621_n_41963

   PIN FE_OFN13687_n_143426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.378 249.792 11.406 ;
      END
   END FE_OFN13687_n_143426

   PIN FE_OFN13692_n_41993
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.834 249.792 6.862 ;
      END
   END FE_OFN13692_n_41993

   PIN FE_OFN14071_n_142964
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.442 0.0 19.47 0.163 ;
      END
   END FE_OFN14071_n_142964

   PIN FE_OFN14164_n_31516
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.234 117.597 69.262 117.76 ;
      END
   END FE_OFN14164_n_31516

   PIN FE_OFN14397_n_140213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.938 0.0 229.966 0.163 ;
      END
   END FE_OFN14397_n_140213

   PIN FE_OFN14901_n_140203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.882 249.792 40.91 ;
      END
   END FE_OFN14901_n_140203

   PIN FE_OFN15072_n_29125
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.754 117.597 208.782 117.76 ;
      END
   END FE_OFN15072_n_29125

   PIN FE_OFN15106_n_30279
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.73 117.597 199.758 117.76 ;
      END
   END FE_OFN15106_n_30279

   PIN FE_OFN15135_n_30145
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 71.282 249.792 71.31 ;
      END
   END FE_OFN15135_n_30145

   PIN FE_OFN15329_n_29953
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 188.274 117.597 188.302 117.76 ;
      END
   END FE_OFN15329_n_29953

   PIN FE_OFN15343_n_30559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 203.634 117.597 203.662 117.76 ;
      END
   END FE_OFN15343_n_30559

   PIN FE_OFN16079_n_41709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.898 0.0 238.926 0.163 ;
      END
   END FE_OFN16079_n_41709

   PIN FE_OFN16087_n_41993
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.666 249.792 55.694 ;
      END
   END FE_OFN16087_n_41993

   PIN FE_OFN16127_n_66979
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.586 0.0 241.614 0.163 ;
      END
   END FE_OFN16127_n_66979

   PIN FE_OFN16313_b_7_6_9
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 244.338 0.0 244.366 0.163 ;
      END
   END FE_OFN16313_b_7_6_9

   PIN FE_OFN17006_n_58282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.466 117.597 124.494 117.76 ;
      END
   END FE_OFN17006_n_58282

   PIN FE_OFN17423_n_8249
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.818 0.0 128.846 0.163 ;
      END
   END FE_OFN17423_n_8249

   PIN FE_OFN17844_n_81895
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 67.762 249.792 67.79 ;
      END
   END FE_OFN17844_n_81895

   PIN FE_OFN17850_n_66751
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 63.666 249.792 63.694 ;
      END
   END FE_OFN17850_n_66751

   PIN FE_OFN17864_n_71795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.042 249.792 29.07 ;
      END
   END FE_OFN17864_n_71795

   PIN FE_OFN17908_n_55576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 2.61 249.792 2.638 ;
      END
   END FE_OFN17908_n_55576

   PIN FE_OFN18784_n_31306
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.538 117.597 111.566 117.76 ;
      END
   END FE_OFN18784_n_31306

   PIN FE_OFN19276_n_28640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.074 117.597 169.102 117.76 ;
      END
   END FE_OFN19276_n_28640

   PIN FE_OFN2321_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.802 117.597 226.83 117.76 ;
      END
   END FE_OFN2321_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_14_

   PIN FE_OFN2322_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 86.834 249.792 86.862 ;
      END
   END FE_OFN2322_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_13_

   PIN FE_OFN4459_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.258 0.0 142.286 0.163 ;
      END
   END FE_OFN4459_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_12_

   PIN FE_OFN4762_n_137230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.738 0.0 18.766 0.082 ;
      END
   END FE_OFN4762_n_137230

   PIN FE_OFN4815_n_143202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.434 0.0 72.462 0.163 ;
      END
   END FE_OFN4815_n_143202

   PIN FE_OFN6162_delay_mul_ln34_unr7_unr8_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 176.818 0.0 176.846 0.163 ;
      END
   END FE_OFN6162_delay_mul_ln34_unr7_unr8_stage2_stallmux_z_13_

   PIN FE_OFN6326_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.762 0.0 139.79 0.163 ;
      END
   END FE_OFN6326_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_7_

   PIN FE_OFN6445_n_64478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 63.09 249.792 63.118 ;
      END
   END FE_OFN6445_n_64478

   PIN FE_OFN6458_n_59534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 242.098 0.0 242.126 0.163 ;
      END
   END FE_OFN6458_n_59534

   PIN FE_OFN6491_n_41960
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 241.266 0.0 241.294 0.163 ;
      END
   END FE_OFN6491_n_41960

   PIN FE_OFN6549_n_41963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.106 249.792 45.134 ;
      END
   END FE_OFN6549_n_41963

   PIN FE_OFN6605_n_140234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.546 0.0 226.574 0.163 ;
      END
   END FE_OFN6605_n_140234

   PIN FE_OFN6626_n_41612
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.37 249.792 48.398 ;
      END
   END FE_OFN6626_n_41612

   PIN FE_OFN6749_n_41995
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 56.306 249.792 56.334 ;
      END
   END FE_OFN6749_n_41995

   PIN FE_OFN6841_n_41015
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.874 249.792 21.902 ;
      END
   END FE_OFN6841_n_41015

   PIN FE_OFN6859_n_143629
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.226 0.0 242.254 0.163 ;
      END
   END FE_OFN6859_n_143629

   PIN FE_OFN8170_n_26637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.082 117.597 132.11 117.76 ;
      END
   END FE_OFN8170_n_26637

   PIN FE_OFN8330_n_31307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.298 117.597 181.326 117.76 ;
      END
   END FE_OFN8330_n_31307

   PIN FE_OFN8366_n_31480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.002 117.597 102.03 117.76 ;
      END
   END FE_OFN8366_n_31480

   PIN FE_OFN8464_n_25371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.578 117.597 230.606 117.76 ;
      END
   END FE_OFN8464_n_25371

   PIN FE_OFN8492_n_29557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 184.37 117.597 184.398 117.76 ;
      END
   END FE_OFN8492_n_29557

   PIN FE_OFN8498_n_28380
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.818 117.597 176.846 117.76 ;
      END
   END FE_OFN8498_n_28380

   PIN FE_OFN8499_n_27857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.002 117.597 142.03 117.76 ;
      END
   END FE_OFN8499_n_27857

   PIN FE_OFN8578_n_29968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 25.138 249.792 25.166 ;
      END
   END FE_OFN8578_n_29968

   PIN FE_OFN8704_n_31118
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.578 249.792 94.606 ;
      END
   END FE_OFN8704_n_31118

   PIN FE_OFN8719_n_25376
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.642 249.792 94.67 ;
      END
   END FE_OFN8719_n_25376

   PIN FE_OFN9239_delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 98.29 249.792 98.318 ;
      END
   END FE_OFN9239_delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_

   PIN FE_OFN9472_b_7_8_8
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 29.426 249.792 29.454 ;
      END
   END FE_OFN9472_b_7_8_8

   PIN FE_OFN9474_b_7_8_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 56.114 249.792 56.142 ;
      END
   END FE_OFN9474_b_7_8_7

   PIN FE_OFN9536_b_7_6_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.818 249.792 32.846 ;
      END
   END FE_OFN9536_b_7_6_15

   PIN FE_OFN9540_b_7_6_14
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 222.962 0.0 222.99 0.163 ;
      END
   END FE_OFN9540_b_7_6_14

   PIN FE_OFN9548_b_7_6_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.026 249.792 7.054 ;
      END
   END FE_OFN9548_b_7_6_11

   PIN FE_OFN9549_b_7_6_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.394 249.792 41.422 ;
      END
   END FE_OFN9549_b_7_6_10

   PIN FE_OFN9558_b_7_6_6
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.066 249.792 22.094 ;
      END
   END FE_OFN9558_b_7_6_6

   PIN FE_OFN9564_b_7_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 56.37 249.792 56.398 ;
      END
   END FE_OFN9564_b_7_6_4

   PIN FE_OFN9577_b_7_6_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 33.33 249.792 33.358 ;
      END
   END FE_OFN9577_b_7_6_1

   PIN FE_OFN9879_b_4_8_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.242 0.0 88.27 0.163 ;
      END
   END FE_OFN9879_b_4_8_3

   PIN delay_mul_ln34_unr4_unr2_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.778 0.0 145.806 0.163 ;
      END
   END delay_mul_ln34_unr4_unr2_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr4_unr2_stage2_stallmux_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.714 0.0 65.742 0.163 ;
      END
   END delay_mul_ln34_unr4_unr2_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr4_unr4_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.01 0.0 113.038 0.163 ;
      END
   END delay_mul_ln34_unr4_unr4_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr4_unr6_stage2_stallmux_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.362 0.0 125.39 0.163 ;
      END
   END delay_mul_ln34_unr4_unr6_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr4_unr6_stage2_stallmux_z_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.546 0.0 114.574 0.163 ;
      END
   END delay_mul_ln34_unr4_unr6_stage2_stallmux_z_8_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.978 249.792 85.006 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr7_unr8_stage2_stallmux_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.098 0.0 154.126 0.163 ;
      END
   END delay_mul_ln34_unr7_unr8_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.906 117.597 145.934 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.122 117.597 139.15 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_q_3_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.93 117.597 218.958 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.066 117.597 142.094 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_4_

   PIN mul_4647_72_n_200
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.018 0.0 4.046 0.163 ;
      END
   END mul_4647_72_n_200

   PIN mul_4647_72_n_224
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.898 0.0 22.926 0.163 ;
      END
   END mul_4647_72_n_224

   PIN mul_4647_72_n_227
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.242 0.0 8.27 0.163 ;
      END
   END mul_4647_72_n_227

   PIN mul_4647_72_n_230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.082 0.0 20.11 0.163 ;
      END
   END mul_4647_72_n_230

   PIN mul_4647_72_n_252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.77 0.0 30.798 0.163 ;
      END
   END mul_4647_72_n_252

   PIN mul_4647_72_n_323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.786 0.0 36.814 0.163 ;
      END
   END mul_4647_72_n_323

   PIN mul_4647_72_n_71
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.378 0.0 11.406 0.163 ;
      END
   END mul_4647_72_n_71

   PIN mul_4649_72_n_77
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.09 0.0 119.118 0.163 ;
      END
   END mul_4649_72_n_77

   PIN mul_4651_72_n_290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.85 0.0 76.878 0.163 ;
      END
   END mul_4651_72_n_290

   PIN mul_4651_72_n_316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.906 0.0 73.934 0.163 ;
      END
   END mul_4651_72_n_316

   PIN mul_4651_72_n_322
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.082 0.0 68.11 0.163 ;
      END
   END mul_4651_72_n_322

   PIN mul_4651_72_n_323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.474 0.0 71.502 0.163 ;
      END
   END mul_4651_72_n_323

   PIN mul_4651_72_n_324
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.154 0.0 71.182 0.163 ;
      END
   END mul_4651_72_n_324

   PIN mul_4664_72_n_213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.994 0.0 27.022 0.163 ;
      END
   END mul_4664_72_n_213

   PIN mul_4664_72_n_214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.93 0.0 66.958 0.163 ;
      END
   END mul_4664_72_n_214

   PIN mul_4664_72_n_285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.082 0.0 36.11 0.163 ;
      END
   END mul_4664_72_n_285

   PIN mul_4664_72_n_55
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.986 0.0 8.014 0.163 ;
      END
   END mul_4664_72_n_55

   PIN mul_4664_72_n_71
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.05 0.0 8.078 0.163 ;
      END
   END mul_4664_72_n_71

   PIN mul_4664_72_n_773
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.674 0.0 34.702 0.163 ;
      END
   END mul_4664_72_n_773

   PIN mul_4698_72_n_117
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 223.474 0.0 223.502 0.163 ;
      END
   END mul_4698_72_n_117

   PIN mul_4700_72_n_53
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.962 249.792 6.99 ;
      END
   END mul_4700_72_n_53

   PIN mul_4700_72_n_69
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 211.314 0.0 211.342 0.163 ;
      END
   END mul_4700_72_n_69

   PIN n_100733
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.89 117.597 195.918 117.76 ;
      END
   END n_100733

   PIN n_100744
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.826 117.597 195.854 117.76 ;
      END
   END n_100744

   PIN n_102607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.81 249.792 29.838 ;
      END
   END n_102607

   PIN n_102890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.746 0.0 149.774 0.163 ;
      END
   END n_102890

   PIN n_103077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.858 117.597 199.886 117.76 ;
      END
   END n_103077

   PIN n_103482
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 86.898 249.792 86.926 ;
      END
   END n_103482

   PIN n_105239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.09 117.597 215.118 117.76 ;
      END
   END n_105239

   PIN n_106473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.954 117.597 195.982 117.76 ;
      END
   END n_106473

   PIN n_107990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.45 0.0 38.478 0.163 ;
      END
   END n_107990

   PIN n_108077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.642 117.597 182.67 117.76 ;
      END
   END n_108077

   PIN n_108091
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.898 249.792 94.926 ;
      END
   END n_108091

   PIN n_108970
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.562 0.0 40.59 0.163 ;
      END
   END n_108970

   PIN n_109766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.57 117.597 203.598 117.76 ;
      END
   END n_109766

   PIN n_110534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.506 117.597 203.534 117.76 ;
      END
   END n_110534

   PIN n_110678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.938 249.792 21.966 ;
      END
   END n_110678

   PIN n_110705
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 114.226 249.792 114.254 ;
      END
   END n_110705

   PIN n_11212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.898 0.0 14.926 0.163 ;
      END
   END n_11212

   PIN n_11214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.314 0.0 115.342 0.163 ;
      END
   END n_11214

   PIN n_114514
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.962 0.0 30.99 0.163 ;
      END
   END n_114514

   PIN n_115085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.386 0.0 30.414 0.163 ;
      END
   END n_115085

   PIN n_115534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.194 117.597 54.222 117.76 ;
      END
   END n_115534

   PIN n_115535
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.13 117.597 46.158 117.76 ;
      END
   END n_115535

   PIN n_115594
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.722 0.0 20.75 0.163 ;
      END
   END n_115594

   PIN n_115658
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.058 0.0 27.086 0.163 ;
      END
   END n_115658

   PIN n_116050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.89 0.0 43.918 0.163 ;
      END
   END n_116050

   PIN n_116051
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.954 0.0 43.982 0.163 ;
      END
   END n_116051

   PIN n_116348
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.978 0.0 37.006 0.163 ;
      END
   END n_116348

   PIN n_116462
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 11.122 0.163 11.15 ;
      END
   END n_116462

   PIN n_116511
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.282 0.0 71.31 0.163 ;
      END
   END n_116511

   PIN n_116767
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.738 0.0 34.766 0.163 ;
      END
   END n_116767

   PIN n_116839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.842 0.0 41.87 0.163 ;
      END
   END n_116839

   PIN n_118700
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.098 0.0 2.126 0.163 ;
      END
   END n_118700

   PIN n_118762
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.25 0.0 19.278 0.163 ;
      END
   END n_118762

   PIN n_118773
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.442 0.163 3.47 ;
      END
   END n_118773

   PIN n_118968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.122 0.0 19.15 0.163 ;
      END
   END n_118968

   PIN n_118969
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.154 0.0 15.182 0.163 ;
      END
   END n_118969

   PIN n_118970
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.282 0.0 15.31 0.163 ;
      END
   END n_118970

   PIN n_119000
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.826 0.0 43.854 0.163 ;
      END
   END n_119000

   PIN n_119073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.506 0.163 75.534 ;
      END
   END n_119073

   PIN n_119481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.482 0.0 18.51 0.163 ;
      END
   END n_119481

   PIN n_119509
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.514 0.0 38.542 0.163 ;
      END
   END n_119509

   PIN n_120297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.162 0.163 10.19 ;
      END
   END n_120297

   PIN n_120453
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.834 0.0 30.862 0.163 ;
      END
   END n_120453

   PIN n_120804
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.306 0.0 48.334 0.163 ;
      END
   END n_120804

   PIN n_120838
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.482 0.163 2.51 ;
      END
   END n_120838

   PIN n_120840
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.93 0.0 18.958 0.163 ;
      END
   END n_120840

   PIN n_121307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.722 0.0 76.75 0.163 ;
      END
   END n_121307

   PIN n_121492
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.898 0.0 30.926 0.163 ;
      END
   END n_121492

   PIN n_121670
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.658 0.0 76.686 0.163 ;
      END
   END n_121670

   PIN n_121988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.242 0.0 16.27 0.163 ;
      END
   END n_121988

   PIN n_122043
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.73 0.163 71.758 ;
      END
   END n_122043

   PIN n_122081
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.93 0.0 26.958 0.163 ;
      END
   END n_122081

   PIN n_122221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.402 0.0 4.43 0.163 ;
      END
   END n_122221

   PIN n_122483
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.242 0.163 56.27 ;
      END
   END n_122483

   PIN n_122484
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.282 0.163 55.31 ;
      END
   END n_122484

   PIN n_122506
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.602 0.163 71.63 ;
      END
   END n_122506

   PIN n_122507
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.842 0.163 25.87 ;
      END
   END n_122507

   PIN n_123326
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.722 0.0 12.75 0.163 ;
      END
   END n_123326

   PIN n_124275
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.53 0.163 52.558 ;
      END
   END n_124275

   PIN n_124317
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.962 0.0 22.99 0.163 ;
      END
   END n_124317

   PIN n_124544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.746 117.597 37.774 117.76 ;
      END
   END n_124544

   PIN n_124640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.066 117.597 46.094 117.76 ;
      END
   END n_124640

   PIN n_124871
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.994 0.0 27.022 0.163 ;
      END
   END n_124871

   PIN n_126137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.618 117.597 37.646 117.76 ;
      END
   END n_126137

   PIN n_127194
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.858 0.0 7.886 0.163 ;
      END
   END n_127194

   PIN n_127226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.386 117.597 38.414 117.76 ;
      END
   END n_127226

   PIN n_127725
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.746 0.163 21.774 ;
      END
   END n_127725

   PIN n_127726
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.162 0.163 18.19 ;
      END
   END n_127726

   PIN n_128154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.858 0.0 7.886 0.163 ;
      END
   END n_128154

   PIN n_128155
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.922 0.0 7.95 0.163 ;
      END
   END n_128155

   PIN n_128174
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.834 0.0 22.862 0.163 ;
      END
   END n_128174

   PIN n_128290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.85 0.163 44.878 ;
      END
   END n_128290

   PIN n_128294
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.522 0.0 9.55 0.163 ;
      END
   END n_128294

   PIN n_129242
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.042 117.597 21.07 117.76 ;
      END
   END n_129242

   PIN n_129244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.698 117.597 27.726 117.76 ;
      END
   END n_129244

   PIN n_129371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.474 117.597 15.502 117.76 ;
      END
   END n_129371

   PIN n_129623
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 99.442 0.163 99.47 ;
      END
   END n_129623

   PIN n_129649
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 84.722 0.163 84.75 ;
      END
   END n_129649

   PIN n_129721
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.21 0.0 4.238 0.163 ;
      END
   END n_129721

   PIN n_130485
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.41 117.597 15.438 117.76 ;
      END
   END n_130485

   PIN n_131556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.498 117.597 32.526 117.76 ;
      END
   END n_131556

   PIN n_133552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.914 0.0 36.942 0.163 ;
      END
   END n_133552

   PIN n_134508
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.186 0.0 19.214 0.163 ;
      END
   END n_134508

   PIN n_135085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.314 0.0 19.342 0.163 ;
      END
   END n_135085

   PIN n_137235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.954 0.0 227.982 0.163 ;
      END
   END n_137235

   PIN n_137837
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.306 0.0 88.334 0.163 ;
      END
   END n_137837

   PIN n_143371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.442 249.792 11.47 ;
      END
   END n_143371

   PIN n_143818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.186 0.0 11.214 0.163 ;
      END
   END n_143818

   PIN n_24537
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 194.738 0.0 194.766 0.163 ;
      END
   END n_24537

   PIN n_24538
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 188.146 0.0 188.174 0.163 ;
      END
   END n_24538

   PIN n_25880
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.074 0.0 169.102 0.163 ;
      END
   END n_25880

   PIN n_25882
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 173.298 0.0 173.326 0.163 ;
      END
   END n_25882

   PIN n_26382
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.97 117.597 145.998 117.76 ;
      END
   END n_26382

   PIN n_26770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.394 117.597 145.422 117.76 ;
      END
   END n_26770

   PIN n_26771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 146.034 117.597 146.062 117.76 ;
      END
   END n_26771

   PIN n_26989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.938 0.0 149.966 0.163 ;
      END
   END n_26989

   PIN n_27355
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 192.114 117.597 192.142 117.76 ;
      END
   END n_27355

   PIN n_28369
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.85 117.597 116.878 117.76 ;
      END
   END n_28369

   PIN n_2842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.866 0.0 10.894 0.163 ;
      END
   END n_2842

   PIN n_28483
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 95.09 249.792 95.118 ;
      END
   END n_28483

   PIN n_28878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.794 117.597 119.822 117.76 ;
      END
   END n_28878

   PIN n_29113
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.962 249.792 94.99 ;
      END
   END n_29113

   PIN n_2937
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.154 0.0 119.182 0.163 ;
      END
   END n_2937

   PIN n_29558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 184.306 117.597 184.334 117.76 ;
      END
   END n_29558

   PIN n_32569
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.218 0.0 47.246 0.163 ;
      END
   END n_32569

   PIN n_32599
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.442 0.0 67.47 0.163 ;
      END
   END n_32599

   PIN n_32677
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.89 0.0 75.918 0.163 ;
      END
   END n_32677

   PIN n_32709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.482 0.0 34.51 0.163 ;
      END
   END n_32709

   PIN n_32886
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.906 0.0 49.934 0.163 ;
      END
   END n_32886

   PIN n_33168
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 25.33 249.792 25.358 ;
      END
   END n_33168

   PIN n_33209
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.042 0.0 93.07 0.163 ;
      END
   END n_33209

   PIN n_33371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 231.922 0.0 231.95 0.163 ;
      END
   END n_33371

   PIN n_34045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.218 0.0 23.246 0.163 ;
      END
   END n_34045

   PIN n_34363
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.266 0.0 81.294 0.163 ;
      END
   END n_34363

   PIN n_34386
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.706 0.0 110.734 0.163 ;
      END
   END n_34386

   PIN n_34739
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.762 249.792 3.79 ;
      END
   END n_34739

   PIN n_35423
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.202 0.0 81.23 0.163 ;
      END
   END n_35423

   PIN n_36289
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.09 0.0 71.118 0.163 ;
      END
   END n_36289

   PIN n_36486
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.938 0.0 93.966 0.163 ;
      END
   END n_36486

   PIN n_36699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.746 0.0 53.774 0.163 ;
      END
   END n_36699

   PIN n_36728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.842 0.0 65.87 0.163 ;
      END
   END n_36728

   PIN n_36741
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.826 249.792 3.854 ;
      END
   END n_36741

   PIN n_36776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.914 0.0 212.942 0.163 ;
      END
   END n_36776

   PIN n_36951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.97 0.0 49.998 0.163 ;
      END
   END n_36951

   PIN n_37371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.002 0.0 46.03 0.163 ;
      END
   END n_37371

   PIN n_37496
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.33 0.0 65.358 0.163 ;
      END
   END n_37496

   PIN n_37823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.786 0.0 76.814 0.163 ;
      END
   END n_37823

   PIN n_38020
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.426 0.0 61.454 0.163 ;
      END
   END n_38020

   PIN n_38377
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.682 0.0 37.71 0.163 ;
      END
   END n_38377

   PIN n_39631
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.618 0.0 37.646 0.163 ;
      END
   END n_39631

   PIN n_40828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.938 0.0 245.966 0.163 ;
      END
   END n_40828

   PIN n_40903
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.066 0.0 70.094 0.163 ;
      END
   END n_40903

   PIN n_43135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.954 249.792 99.982 ;
      END
   END n_43135

   PIN n_43460
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 69.106 249.792 69.134 ;
      END
   END n_43460

   PIN n_43886
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.842 249.792 33.87 ;
      END
   END n_43886

   PIN n_43887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.586 249.792 33.614 ;
      END
   END n_43887

   PIN n_43927
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 76.786 249.792 76.814 ;
      END
   END n_43927

   PIN n_43959
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.826 249.792 11.854 ;
      END
   END n_43959

   PIN n_44225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.45 249.792 70.478 ;
      END
   END n_44225

   PIN n_44595
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 100.018 249.792 100.046 ;
      END
   END n_44595

   PIN n_44641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.89 249.792 3.918 ;
      END
   END n_44641

   PIN n_44714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.73 249.792 55.758 ;
      END
   END n_44714

   PIN n_44715
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 56.178 249.792 56.206 ;
      END
   END n_44715

   PIN n_44776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 36.594 249.792 36.622 ;
      END
   END n_44776

   PIN n_44777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 36.658 249.792 36.686 ;
      END
   END n_44777

   PIN n_45142
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.594 249.792 44.622 ;
      END
   END n_45142

   PIN n_45217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 79.218 249.792 79.246 ;
      END
   END n_45217

   PIN n_45222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.546 0.0 130.574 0.163 ;
      END
   END n_45222

   PIN n_45299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 184.306 0.0 184.334 0.163 ;
      END
   END n_45299

   PIN n_45510
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.498 0.0 112.526 0.163 ;
      END
   END n_45510

   PIN n_45631
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.402 0.0 84.43 0.163 ;
      END
   END n_45631

   PIN n_45632
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.242 0.0 80.27 0.163 ;
      END
   END n_45632

   PIN n_45699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 2.674 249.792 2.702 ;
      END
   END n_45699

   PIN n_45883
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 76.722 249.792 76.75 ;
      END
   END n_45883

   PIN n_46067
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.61 0.0 130.638 0.163 ;
      END
   END n_46067

   PIN n_46081
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.21 249.792 52.238 ;
      END
   END n_46081

   PIN n_46203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 172.914 0.0 172.942 0.163 ;
      END
   END n_46203

   PIN n_46332
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.498 249.792 48.526 ;
      END
   END n_46332

   PIN n_46335
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 4.082 249.792 4.11 ;
      END
   END n_46335

   PIN n_46361
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.69 249.792 32.718 ;
      END
   END n_46361

   PIN n_46369
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.594 249.792 84.622 ;
      END
   END n_46369

   PIN n_46370
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.402 249.792 84.43 ;
      END
   END n_46370

   PIN n_46467
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 60.338 249.792 60.366 ;
      END
   END n_46467

   PIN n_46468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 60.402 249.792 60.43 ;
      END
   END n_46468

   PIN n_46540
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.146 249.792 52.174 ;
      END
   END n_46540

   PIN n_46576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.242 0.0 112.27 0.163 ;
      END
   END n_46576

   PIN n_46582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 63.794 249.792 63.822 ;
      END
   END n_46582

   PIN n_46583
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 2.738 249.792 2.766 ;
      END
   END n_46583

   PIN n_46659
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.89 249.792 11.918 ;
      END
   END n_46659

   PIN n_46661
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.514 0.0 110.542 0.163 ;
      END
   END n_46661

   PIN n_46668
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.754 249.792 48.782 ;
      END
   END n_46668

   PIN n_46669
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.402 249.792 44.43 ;
      END
   END n_46669

   PIN n_46676
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 238.194 0.0 238.222 0.163 ;
      END
   END n_46676

   PIN n_46872
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.002 249.792 22.03 ;
      END
   END n_46872

   PIN n_46916
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.834 0.0 94.862 0.163 ;
      END
   END n_46916

   PIN n_46917
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.642 0.0 86.67 0.163 ;
      END
   END n_46917

   PIN n_47149
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.042 249.792 37.07 ;
      END
   END n_47149

   PIN n_47248
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 79.346 249.792 79.374 ;
      END
   END n_47248

   PIN n_47260
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.226 0.0 138.254 0.163 ;
      END
   END n_47260

   PIN n_47323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.498 0.0 216.526 0.163 ;
      END
   END n_47323

   PIN n_47423
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.53 249.792 84.558 ;
      END
   END n_47423

   PIN n_47856
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.938 0.0 53.966 0.163 ;
      END
   END n_47856

   PIN n_47857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.922 0.0 63.95 0.163 ;
      END
   END n_47857

   PIN n_49211
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.194 0.0 38.222 0.163 ;
      END
   END n_49211

   PIN n_49947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.106 249.792 29.134 ;
      END
   END n_49947

   PIN n_50245
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 86.77 249.792 86.798 ;
      END
   END n_50245

   PIN n_50316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.578 249.792 110.606 ;
      END
   END n_50316

   PIN n_50589
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 71.346 249.792 71.374 ;
      END
   END n_50589

   PIN n_50941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.002 0.0 246.03 0.163 ;
      END
   END n_50941

   PIN n_51049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.514 0.0 134.542 0.163 ;
      END
   END n_51049

   PIN n_51080
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 188.21 0.0 188.238 0.163 ;
      END
   END n_51080

   PIN n_51152
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.234 0.0 109.262 0.163 ;
      END
   END n_51152

   PIN n_51247
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.658 249.792 44.686 ;
      END
   END n_51247

   PIN n_52208
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.354 249.792 26.382 ;
      END
   END n_52208

   PIN n_52412
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 63.154 249.792 63.182 ;
      END
   END n_52412

   PIN n_52666
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 59.89 249.792 59.918 ;
      END
   END n_52666

   PIN n_52803
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.466 249.792 84.494 ;
      END
   END n_52803

   PIN n_52852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.386 249.792 102.414 ;
      END
   END n_52852

   PIN n_53092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.162 0.0 138.19 0.163 ;
      END
   END n_53092

   PIN n_53255
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 87.026 249.792 87.054 ;
      END
   END n_53255

   PIN n_53257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 222.066 0.0 222.094 0.163 ;
      END
   END n_53257

   PIN n_53297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 67.826 249.792 67.854 ;
      END
   END n_53297

   PIN n_53524
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.106 249.792 37.134 ;
      END
   END n_53524

   PIN n_53555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 98.354 249.792 98.382 ;
      END
   END n_53555

   PIN n_53566
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.482 249.792 106.51 ;
      END
   END n_53566

   PIN n_53983
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.65 0.0 81.678 0.163 ;
      END
   END n_53983

   PIN n_53996
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.594 249.792 52.622 ;
      END
   END n_53996

   PIN n_54311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.298 0.0 61.326 0.163 ;
      END
   END n_54311

   PIN n_54338
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.17 249.792 77.198 ;
      END
   END n_54338

   PIN n_54688
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 17.458 249.792 17.486 ;
      END
   END n_54688

   PIN n_54944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.314 117.597 139.342 117.76 ;
      END
   END n_54944

   PIN n_54954
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.25 117.597 115.278 117.76 ;
      END
   END n_54954

   PIN n_54986
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.642 249.792 110.67 ;
      END
   END n_54986

   PIN n_55042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.402 249.792 92.43 ;
      END
   END n_55042

   PIN n_55157
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.258 117.597 158.286 117.76 ;
      END
   END n_55157

   PIN n_55513
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 17.586 249.792 17.614 ;
      END
   END n_55513

   PIN n_5555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 6.386 249.792 6.414 ;
      END
   END n_5555

   PIN n_55597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.01 249.792 41.038 ;
      END
   END n_55597

   PIN n_55598
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.17 249.792 29.198 ;
      END
   END n_55598

   PIN n_55674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 184.434 0.0 184.462 0.163 ;
      END
   END n_55674

   PIN n_55702
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.594 0.0 100.622 0.163 ;
      END
   END n_55702

   PIN n_55723
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.05 0.0 120.078 0.163 ;
      END
   END n_55723

   PIN n_55740
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.97 0.0 145.998 0.163 ;
      END
   END n_55740

   PIN n_55766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.97 249.792 33.998 ;
      END
   END n_55766

   PIN n_56659
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.794 249.792 55.822 ;
      END
   END n_56659

   PIN n_56808
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.018 249.792 92.046 ;
      END
   END n_56808

   PIN n_56899
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.658 249.792 84.686 ;
      END
   END n_56899

   PIN n_57040
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.626 0.0 80.654 0.163 ;
      END
   END n_57040

   PIN n_57135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.426 0.163 29.454 ;
      END
   END n_57135

   PIN n_57460
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.842 0.0 137.87 0.163 ;
      END
   END n_57460

   PIN n_57673
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 179.634 0.0 179.662 0.163 ;
      END
   END n_57673

   PIN n_57704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.034 0.0 242.062 0.163 ;
      END
   END n_57704

   PIN n_57712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.266 0.0 161.294 0.163 ;
      END
   END n_57712

   PIN n_57713
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.674 0.0 162.702 0.163 ;
      END
   END n_57713

   PIN n_57714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.442 0.0 163.47 0.163 ;
      END
   END n_57714

   PIN n_57823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 37.81 249.792 37.838 ;
      END
   END n_57823

   PIN n_57902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.346 117.597 111.374 117.76 ;
      END
   END n_57902

   PIN n_57982
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 153.714 117.597 153.742 117.76 ;
      END
   END n_57982

   PIN n_58071
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.282 0.0 239.31 0.163 ;
      END
   END n_58071

   PIN n_58207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.098 0.0 242.126 0.163 ;
      END
   END n_58207

   PIN n_58229
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.698 249.792 99.726 ;
      END
   END n_58229

   PIN n_58234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 106.098 249.792 106.126 ;
      END
   END n_58234

   PIN n_58257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.034 117.597 162.062 117.76 ;
      END
   END n_58257

   PIN n_58264
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.554 117.597 133.582 117.76 ;
      END
   END n_58264

   PIN n_58283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.77 117.597 126.798 117.76 ;
      END
   END n_58283

   PIN n_58292
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.29 0.0 138.318 0.163 ;
      END
   END n_58292

   PIN n_58507
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.346 0.0 247.374 0.163 ;
      END
   END n_58507

   PIN n_59057
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.074 117.597 153.102 117.76 ;
      END
   END n_59057

   PIN n_59287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.586 117.597 161.614 117.76 ;
      END
   END n_59287

   PIN n_59495
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.586 0.0 153.614 0.163 ;
      END
   END n_59495

   PIN n_59615
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.546 249.792 106.574 ;
      END
   END n_59615

   PIN n_59894
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.218 0.0 15.246 0.163 ;
      END
   END n_59894

   PIN n_60087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.514 249.792 110.542 ;
      END
   END n_60087

   PIN n_60088
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 134.514 117.597 134.542 117.76 ;
      END
   END n_60088

   PIN n_60104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 47.602 249.792 47.63 ;
      END
   END n_60104

   PIN n_60139
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.082 249.792 92.11 ;
      END
   END n_60139

   PIN n_60261
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.146 249.792 92.174 ;
      END
   END n_60261

   PIN n_60264
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.962 117.597 158.99 117.76 ;
      END
   END n_60264

   PIN n_60317
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.066 117.597 126.094 117.76 ;
      END
   END n_60317

   PIN n_60318
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.002 117.597 126.03 117.76 ;
      END
   END n_60318

   PIN n_60377
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.002 249.792 70.03 ;
      END
   END n_60377

   PIN n_60444
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.45 249.792 102.478 ;
      END
   END n_60444

   PIN n_60543
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.434 249.792 48.462 ;
      END
   END n_60543

   PIN n_60569
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.754 0.0 176.782 0.163 ;
      END
   END n_60569

   PIN n_60575
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.122 0.0 163.15 0.163 ;
      END
   END n_60575

   PIN n_60581
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.69 0.0 176.718 0.163 ;
      END
   END n_60581

   PIN n_60661
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.074 117.597 113.102 117.76 ;
      END
   END n_60661

   PIN n_60763
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.074 249.792 33.102 ;
      END
   END n_60763

   PIN n_60770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.074 117.597 137.102 117.76 ;
      END
   END n_60770

   PIN n_61110
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.53 117.597 84.558 117.76 ;
      END
   END n_61110

   PIN n_61151
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.306 0.0 112.334 0.163 ;
      END
   END n_61151

   PIN n_61597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.898 249.792 6.926 ;
      END
   END n_61597

   PIN n_61600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.666 249.792 47.694 ;
      END
   END n_61600

   PIN n_61622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.714 0.0 153.742 0.163 ;
      END
   END n_61622

   PIN n_61766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.65 0.0 89.678 0.163 ;
      END
   END n_61766

   PIN n_61876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.818 117.597 160.846 117.76 ;
      END
   END n_61876

   PIN n_61877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.754 117.597 160.782 117.76 ;
      END
   END n_61877

   PIN n_61881
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 157.554 117.597 157.582 117.76 ;
      END
   END n_61881

   PIN n_61896
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.458 117.597 129.486 117.76 ;
      END
   END n_61896

   PIN n_62357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.594 117.597 84.622 117.76 ;
      END
   END n_62357

   PIN n_62360
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.194 249.792 14.222 ;
      END
   END n_62360

   PIN n_62401
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.33 0.0 105.358 0.163 ;
      END
   END n_62401

   PIN n_62504
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.066 0.0 246.094 0.163 ;
      END
   END n_62504

   PIN n_62647
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.082 0.0 164.11 0.163 ;
      END
   END n_62647

   PIN n_62807
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.394 117.597 65.422 117.76 ;
      END
   END n_62807

   PIN n_62808
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.41 117.597 71.438 117.76 ;
      END
   END n_62808

   PIN n_62998
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.986 117.597 96.014 117.76 ;
      END
   END n_62998

   PIN n_63006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 34.034 249.792 34.062 ;
      END
   END n_63006

   PIN n_63048
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 71.41 249.792 71.438 ;
      END
   END n_63048

   PIN n_63049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.514 249.792 70.542 ;
      END
   END n_63049

   PIN n_63050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.378 0.0 155.406 0.163 ;
      END
   END n_63050

   PIN n_63051
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.146 0.0 148.174 0.163 ;
      END
   END n_63051

   PIN n_63137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 17.714 249.792 17.742 ;
      END
   END n_63137

   PIN n_63203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 234.29 0.0 234.318 0.163 ;
      END
   END n_63203

   PIN n_63244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.202 117.597 161.23 117.76 ;
      END
   END n_63244

   PIN n_63246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.01 117.597 169.038 117.76 ;
      END
   END n_63246

   PIN n_63253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 189.618 117.597 189.646 117.76 ;
      END
   END n_63253

   PIN n_63258
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.25 117.597 211.278 117.76 ;
      END
   END n_63258

   PIN n_63272
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.642 0.0 182.67 0.163 ;
      END
   END n_63272

   PIN n_63359
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 185.074 0.0 185.102 0.163 ;
      END
   END n_63359

   PIN n_63530
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.458 117.597 153.486 117.76 ;
      END
   END n_63530

   PIN n_63531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.042 117.597 157.07 117.76 ;
      END
   END n_63531

   PIN n_63563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 86.962 249.792 86.99 ;
      END
   END n_63563

   PIN n_6357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.394 0.0 121.422 0.163 ;
      END
   END n_6357

   PIN n_63724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.258 249.792 14.286 ;
      END
   END n_63724

   PIN n_64400
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.794 0.0 103.822 0.163 ;
      END
   END n_64400

   PIN n_64412
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.618 0.0 149.646 0.163 ;
      END
   END n_64412

   PIN n_64413
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.85 0.0 148.878 0.163 ;
      END
   END n_64413

   PIN n_64467
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.762 117.597 99.79 117.76 ;
      END
   END n_64467

   PIN n_64527
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 63.73 249.792 63.758 ;
      END
   END n_64527

   PIN n_64551
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.138 117.597 169.166 117.76 ;
      END
   END n_64551

   PIN n_64555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.778 117.597 145.806 117.76 ;
      END
   END n_64555

   PIN n_64556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.194 117.597 142.222 117.76 ;
      END
   END n_64556

   PIN n_64558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.818 117.597 128.846 117.76 ;
      END
   END n_64558

   PIN n_64834
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.354 0.0 138.382 0.163 ;
      END
   END n_64834

   PIN n_64921
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.906 249.792 33.934 ;
      END
   END n_64921

   PIN n_64944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.386 249.792 70.414 ;
      END
   END n_64944

   PIN n_64988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.506 0.0 91.534 0.163 ;
      END
   END n_64988

   PIN n_65021
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.282 117.597 159.31 117.76 ;
      END
   END n_65021

   PIN n_65147
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.946 117.597 152.974 117.76 ;
      END
   END n_65147

   PIN n_65154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 13.938 249.792 13.966 ;
      END
   END n_65154

   PIN n_65353
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.898 117.597 142.926 117.76 ;
      END
   END n_65353

   PIN n_65402
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 184.434 0.0 184.462 0.163 ;
      END
   END n_65402

   PIN n_65488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.178 249.792 48.206 ;
      END
   END n_65488

   PIN n_65500
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 153.65 117.597 153.678 117.76 ;
      END
   END n_65500

   PIN n_65528
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 184.37 0.0 184.398 0.163 ;
      END
   END n_65528

   PIN n_65632
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.186 117.597 155.214 117.76 ;
      END
   END n_65632

   PIN n_65654
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.522 117.597 153.55 117.76 ;
      END
   END n_65654

   PIN n_65680
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.65 0.0 153.678 0.163 ;
      END
   END n_65680

   PIN n_65751
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.266 117.597 153.294 117.76 ;
      END
   END n_65751

   PIN n_65798
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.154 117.597 95.182 117.76 ;
      END
   END n_65798

   PIN n_65952
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.114 0.0 128.142 0.163 ;
      END
   END n_65952

   PIN n_65974
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.506 249.792 11.534 ;
      END
   END n_65974

   PIN n_66586
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 11.186 249.792 11.214 ;
      END
   END n_66586

   PIN n_66611
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 142.13 0.0 142.158 0.163 ;
      END
   END n_66611

   PIN n_66722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.154 117.597 215.182 117.76 ;
      END
   END n_66722

   PIN n_66841
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.042 249.792 77.07 ;
      END
   END n_66841

   PIN n_67151
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.122 117.597 155.15 117.76 ;
      END
   END n_67151

   PIN n_67191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.13 117.597 142.158 117.76 ;
      END
   END n_67191

   PIN n_71276
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 26.034 249.792 26.062 ;
      END
   END n_71276

   PIN n_71277
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.874 249.792 29.902 ;
      END
   END n_71277

   PIN n_71278
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 25.394 249.792 25.422 ;
      END
   END n_71278

   PIN n_71434
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 25.97 249.792 25.998 ;
      END
   END n_71434

   PIN n_71435
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.418 249.792 26.446 ;
      END
   END n_71435

   PIN n_71444
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.666 0.0 103.694 0.163 ;
      END
   END n_71444

   PIN n_71763
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.17 249.792 37.198 ;
      END
   END n_71763

   PIN n_71770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 75.506 249.792 75.534 ;
      END
   END n_71770

   PIN n_72006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.914 117.597 148.942 117.76 ;
      END
   END n_72006

   PIN n_72275
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.234 249.792 77.262 ;
      END
   END n_72275

   PIN n_77145
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.058 117.597 155.086 117.76 ;
      END
   END n_77145

   PIN n_77670
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.642 249.792 6.67 ;
      END
   END n_77670

   PIN n_77995
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.082 117.597 196.11 117.76 ;
      END
   END n_77995

   PIN n_78280
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 76.85 249.792 76.878 ;
      END
   END n_78280

   PIN n_78473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.53 117.597 140.558 117.76 ;
      END
   END n_78473

   PIN n_8031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.738 0.0 10.766 0.163 ;
      END
   END n_8031

   PIN n_82565
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 70.002 249.792 70.03 ;
      END
   END n_82565

   PIN n_83303
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 87.026 249.792 87.054 ;
      END
   END n_83303

   PIN n_8403
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.666 0.0 23.694 0.163 ;
      END
   END n_8403

   PIN n_84678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.298 249.792 77.326 ;
      END
   END n_84678

   PIN n_85584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.442 0.0 131.47 0.163 ;
      END
   END n_85584

   PIN n_88925
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 95.986 249.792 96.014 ;
      END
   END n_88925

   PIN n_91246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 87.09 249.792 87.118 ;
      END
   END n_91246

   PIN n_91249
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.61 249.792 106.638 ;
      END
   END n_91249

   PIN n_91279
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.21 249.792 92.238 ;
      END
   END n_91279

   PIN n_91722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.858 249.792 55.886 ;
      END
   END n_91722

   PIN n_91724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.61 117.597 106.638 117.76 ;
      END
   END n_91724

   PIN n_92857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 60.082 249.792 60.11 ;
      END
   END n_92857

   PIN n_94960
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 95.026 249.792 95.054 ;
      END
   END n_94960

   PIN n_96293
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.626 117.597 136.654 117.76 ;
      END
   END n_96293

   PIN n_97165
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 87.154 249.792 87.182 ;
      END
   END n_97165

   PIN n_97291
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.746 0.0 61.774 0.163 ;
      END
   END n_97291

   PIN FE_OFN10008_b_4_4_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.354 0.0 42.382 0.163 ;
      END
   END FE_OFN10008_b_4_4_11

   PIN FE_OFN10010_b_4_4_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.418 0.0 42.446 0.163 ;
      END
   END FE_OFN10010_b_4_4_10

   PIN FE_OFN10012_b_4_4_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.37 0.0 48.398 0.163 ;
      END
   END FE_OFN10012_b_4_4_9

   PIN FE_OFN10014_b_4_4_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.834 0.0 14.862 0.163 ;
      END
   END FE_OFN10014_b_4_4_8

   PIN FE_OFN10015_b_4_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.386 0.0 38.414 0.163 ;
      END
   END FE_OFN10015_b_4_4_7

   PIN FE_OFN10022_b_4_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.546 0.0 34.574 0.163 ;
      END
   END FE_OFN10022_b_4_4_5

   PIN FE_OFN10023_b_4_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.954 0.0 35.982 0.163 ;
      END
   END FE_OFN10023_b_4_4_5

   PIN FE_OFN10027_b_4_4_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.922 0.0 31.95 0.163 ;
      END
   END FE_OFN10027_b_4_4_3

   PIN FE_OFN10031_b_4_4_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.314 0.0 51.342 0.163 ;
      END
   END FE_OFN10031_b_4_4_2

   PIN FE_OFN10037_b_4_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.914 0.0 20.942 0.163 ;
      END
   END FE_OFN10037_b_4_4_0

   PIN FE_OFN10082_b_4_2_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.41 0.0 47.438 0.163 ;
      END
   END FE_OFN10082_b_4_2_12

   PIN FE_OFN10084_b_4_2_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.746 0.0 53.774 0.163 ;
      END
   END FE_OFN10084_b_4_2_11

   PIN FE_OFN10086_b_4_2_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 57.586 0.0 57.614 0.163 ;
      END
   END FE_OFN10086_b_4_2_10

   PIN FE_OFN10088_b_4_2_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.842 0.0 49.87 0.163 ;
      END
   END FE_OFN10088_b_4_2_9

   PIN FE_OFN10090_b_4_2_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.706 0.0 30.734 0.163 ;
      END
   END FE_OFN10090_b_4_2_8

   PIN FE_OFN10093_b_4_2_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.186 0.0 19.214 0.163 ;
      END
   END FE_OFN10093_b_4_2_7

   PIN FE_OFN10098_b_4_2_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.082 0.0 28.11 0.082 ;
      END
   END FE_OFN10098_b_4_2_5

   PIN FE_OFN10100_b_4_2_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.866 0.0 18.894 0.082 ;
      END
   END FE_OFN10100_b_4_2_4

   PIN FE_OFN10102_b_4_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 49.906 0.0 49.934 0.082 ;
      END
   END FE_OFN10102_b_4_2_3

   PIN FE_OFN10104_b_4_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 57.202 0.0 57.23 0.163 ;
      END
   END FE_OFN10104_b_4_2_2

   PIN FE_OFN10105_b_4_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.874 0.0 53.902 0.163 ;
      END
   END FE_OFN10105_b_4_2_2

   PIN FE_OFN10106_b_4_2_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.322 0.0 38.35 0.163 ;
      END
   END FE_OFN10106_b_4_2_1

   PIN FE_OFN10110_b_4_2_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.162 0.0 58.19 0.082 ;
      END
   END FE_OFN10110_b_4_2_0

   PIN FE_OFN11414_n_140210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.41 0.0 191.438 0.163 ;
      END
   END FE_OFN11414_n_140210

   PIN FE_OFN11419_n_140210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.71 18.29 249.792 18.318 ;
      END
   END FE_OFN11419_n_140210

   PIN FE_OFN11481_n_140205
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 9.65 249.792 9.678 ;
      END
   END FE_OFN11481_n_140205

   PIN FE_OFN11522_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 2.546 249.792 2.574 ;
      END
   END FE_OFN11522_n_140234

   PIN FE_OFN11557_n_137230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.618 0.0 53.646 0.163 ;
      END
   END FE_OFN11557_n_137230

   PIN FE_OFN11558_n_137230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.642 0.0 22.67 0.163 ;
      END
   END FE_OFN11558_n_137230

   PIN FE_OFN11607_n_39244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.386 0.0 70.414 0.163 ;
      END
   END FE_OFN11607_n_39244

   PIN FE_OFN11703_n_36821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.682 0.0 53.71 0.163 ;
      END
   END FE_OFN11703_n_36821

   PIN FE_OFN11879_n_143202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.474 0.0 71.502 0.163 ;
      END
   END FE_OFN11879_n_143202

   PIN FE_OFN11932_n_142850
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.05 0.0 96.078 0.163 ;
      END
   END FE_OFN11932_n_142850

   PIN FE_OFN12024_n_41611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.954 249.792 11.982 ;
      END
   END FE_OFN12024_n_41611

   PIN FE_OFN12028_n_143507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.458 0.0 73.486 0.163 ;
      END
   END FE_OFN12028_n_143507

   PIN FE_OFN12037_n_143629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.41 0.0 247.438 0.163 ;
      END
   END FE_OFN12037_n_143629

   PIN FE_OFN12040_n_143629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.642 0.0 246.67 0.163 ;
      END
   END FE_OFN12040_n_143629

   PIN FE_OFN12061_n_143423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.538 249.792 55.566 ;
      END
   END FE_OFN12061_n_143423

   PIN FE_OFN12085_n_143619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.922 0.0 95.95 0.163 ;
      END
   END FE_OFN12085_n_143619

   PIN FE_OFN12624_n_143670
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 36.914 249.792 36.942 ;
      END
   END FE_OFN12624_n_143670

   PIN FE_OFN12632_n_143496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.77 249.792 6.798 ;
      END
   END FE_OFN12632_n_143496

   PIN FE_OFN12753_n_142961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.098 0.0 50.126 0.163 ;
      END
   END FE_OFN12753_n_142961

   PIN FE_OFN12761_n_41012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 28.978 249.792 29.006 ;
      END
   END FE_OFN12761_n_41012

   PIN FE_OFN12764_n_41015
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.434 249.792 40.462 ;
      END
   END FE_OFN12764_n_41015

   PIN FE_OFN12968_n_112030
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.65 0.0 49.678 0.163 ;
      END
   END FE_OFN12968_n_112030

   PIN FE_OFN13044_n_40829
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 36.85 249.792 36.878 ;
      END
   END FE_OFN13044_n_40829

   PIN FE_OFN13226_n_143481
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 29.362 249.792 29.39 ;
      END
   END FE_OFN13226_n_143481

   PIN FE_OFN13233_n_143479
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.858 0.0 231.886 0.163 ;
      END
   END FE_OFN13233_n_143479

   PIN FE_OFN13239_n_41374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 15.346 249.792 15.374 ;
      END
   END FE_OFN13239_n_41374

   PIN FE_OFN13242_n_41374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.754 249.792 32.782 ;
      END
   END FE_OFN13242_n_41374

   PIN FE_OFN13246_n_143370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.282 0.0 247.31 0.163 ;
      END
   END FE_OFN13246_n_143370

   PIN FE_OFN13253_n_143369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.818 249.792 40.846 ;
      END
   END FE_OFN13253_n_143369

   PIN FE_OFN13297_n_143032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.322 0.0 70.35 0.163 ;
      END
   END FE_OFN13297_n_143032

   PIN FE_OFN13347_n_142796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.13 0.0 38.158 0.163 ;
      END
   END FE_OFN13347_n_142796

   PIN FE_OFN13348_n_142796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.738 0.0 66.766 0.163 ;
      END
   END FE_OFN13348_n_142796

   PIN FE_OFN13393_n_41612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.306 249.792 48.334 ;
      END
   END FE_OFN13393_n_41612

   PIN FE_OFN13450_n_41900
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.53 249.792 52.558 ;
      END
   END FE_OFN13450_n_41900

   PIN FE_OFN13460_n_42034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.818 249.792 48.846 ;
      END
   END FE_OFN13460_n_42034

   PIN FE_OFN13515_n_112357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.77 0.0 30.798 0.163 ;
      END
   END FE_OFN13515_n_112357

   PIN FE_OFN13525_n_137232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.778 0.0 49.806 0.163 ;
      END
   END FE_OFN13525_n_137232

   PIN FE_OFN13528_n_137233
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.13 249.792 14.158 ;
      END
   END FE_OFN13528_n_137233

   PIN FE_OFN13529_n_137233
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.29 249.792 26.318 ;
      END
   END FE_OFN13529_n_137233

   PIN FE_OFN13672_n_143509
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.338 0.0 52.366 0.163 ;
      END
   END FE_OFN13672_n_143509

   PIN FE_OFN13686_n_143426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 247.73 0.0 247.758 0.163 ;
      END
   END FE_OFN13686_n_143426

   PIN FE_OFN13777_n_41686
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.65 0.0 57.678 0.163 ;
      END
   END FE_OFN13777_n_41686

   PIN FE_OFN13787_n_41960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.09 249.792 7.118 ;
      END
   END FE_OFN13787_n_41960

   PIN FE_OFN13789_n_41995
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 13.682 249.792 13.71 ;
      END
   END FE_OFN13789_n_41995

   PIN FE_OFN13796_n_41995
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.778 249.792 33.806 ;
      END
   END FE_OFN13796_n_41995

   PIN FE_OFN13864_n_41964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 37.746 249.792 37.774 ;
      END
   END FE_OFN13864_n_41964

   PIN FE_OFN14082_n_142962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.626 0.0 64.654 0.163 ;
      END
   END FE_OFN14082_n_142962

   PIN FE_OFN14361_n_143300
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.13 0.0 78.158 0.082 ;
      END
   END FE_OFN14361_n_143300

   PIN FE_OFN14401_n_142794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.098 0.0 90.126 0.163 ;
      END
   END FE_OFN14401_n_142794

   PIN FE_OFN14406_n_31761
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.362 0.0 61.39 0.163 ;
      END
   END FE_OFN14406_n_31761

   PIN FE_OFN14899_n_140203
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.73 0.0 247.758 0.163 ;
      END
   END FE_OFN14899_n_140203

   PIN FE_OFN15134_n_30145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 63.026 249.792 63.054 ;
      END
   END FE_OFN15134_n_30145

   PIN FE_OFN15168_n_31480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.034 249.792 106.062 ;
      END
   END FE_OFN15168_n_31480

   PIN FE_OFN15328_n_29953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.45 0.0 230.478 0.163 ;
      END
   END FE_OFN15328_n_29953

   PIN FE_OFN15342_n_30559
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 230.45 0.0 230.478 0.163 ;
      END
   END FE_OFN15342_n_30559

   PIN FE_OFN16113_n_42033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 228.018 0.0 228.046 0.163 ;
      END
   END FE_OFN16113_n_42033

   PIN FE_OFN17005_n_58282
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.738 117.597 226.766 117.76 ;
      END
   END FE_OFN17005_n_58282

   PIN FE_OFN17026_n_66756
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 102.386 249.792 102.414 ;
      END
   END FE_OFN17026_n_66756

   PIN FE_OFN17099_n_53555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 106.482 249.792 106.51 ;
      END
   END FE_OFN17099_n_53555

   PIN FE_OFN17825_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.914 249.792 84.942 ;
      END
   END FE_OFN17825_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_12_

   PIN FE_OFN17835_n_84330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.154 0.0 247.182 0.163 ;
      END
   END FE_OFN17835_n_84330

   PIN FE_OFN17869_n_65432
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.218 0.0 247.246 0.163 ;
      END
   END FE_OFN17869_n_65432

   PIN FE_OFN17921_n_57488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 3.506 249.792 3.534 ;
      END
   END FE_OFN17921_n_57488

   PIN FE_OFN17931_n_41611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.642 0.0 238.67 0.163 ;
      END
   END FE_OFN17931_n_41611

   PIN FE_OFN18301_b_4_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.25 0.0 51.278 0.163 ;
      END
   END FE_OFN18301_b_4_4_4

   PIN FE_OFN18306_b_4_8_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.562 0.0 80.59 0.163 ;
      END
   END FE_OFN18306_b_4_8_5

   PIN FE_OFN18401_n_31516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 60.018 249.792 60.046 ;
      END
   END FE_OFN18401_n_31516

   PIN FE_OFN18434_n_27857
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.066 0.0 238.094 0.163 ;
      END
   END FE_OFN18434_n_27857

   PIN FE_OFN18783_n_31306
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.602 0.0 111.63 0.163 ;
      END
   END FE_OFN18783_n_31306

   PIN FE_OFN18962_n_41993
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.25 249.792 11.278 ;
      END
   END FE_OFN18962_n_41993

   PIN FE_OFN18995_n_41993
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 242.162 0.0 242.19 0.163 ;
      END
   END FE_OFN18995_n_41993

   PIN FE_OFN2320_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.842 117.597 241.87 117.76 ;
      END
   END FE_OFN2320_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_14_

   PIN FE_OFN4455_n_10397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.458 0.0 57.486 0.163 ;
      END
   END FE_OFN4455_n_10397

   PIN FE_OFN4458_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 142.322 0.0 142.35 0.163 ;
      END
   END FE_OFN4458_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_12_

   PIN FE_OFN4574_n_142961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.018 0.0 36.046 0.163 ;
      END
   END FE_OFN4574_n_142961

   PIN FE_OFN4623_n_142793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 49.778 0.0 49.806 0.082 ;
      END
   END FE_OFN4623_n_142793

   PIN FE_OFN4667_n_137232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.338 0.0 28.366 0.163 ;
      END
   END FE_OFN4667_n_137232

   PIN FE_OFN4683_n_143620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.962 0.0 78.99 0.163 ;
      END
   END FE_OFN4683_n_143620

   PIN FE_OFN4730_n_143033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.994 0.0 83.022 0.163 ;
      END
   END FE_OFN4730_n_143033

   PIN FE_OFN4781_n_143003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.898 0.0 38.926 0.163 ;
      END
   END FE_OFN4781_n_143003

   PIN FE_OFN4821_n_143199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.89 0.0 35.918 0.163 ;
      END
   END FE_OFN4821_n_143199

   PIN FE_OFN4837_n_140222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.25 0.0 51.278 0.163 ;
      END
   END FE_OFN4837_n_140222

   PIN FE_OFN4869_n_143507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.858 0.0 31.886 0.163 ;
      END
   END FE_OFN4869_n_143507

   PIN FE_OFN4891_n_140207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.81 0.0 53.838 0.163 ;
      END
   END FE_OFN4891_n_140207

   PIN FE_OFN6426_n_45151
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.722 249.792 52.75 ;
      END
   END FE_OFN6426_n_45151

   PIN FE_OFN6603_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 48.626 249.792 48.654 ;
      END
   END FE_OFN6603_n_140234

   PIN FE_OFN6604_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.71 40.562 249.792 40.59 ;
      END
   END FE_OFN6604_n_140234

   PIN FE_OFN6610_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.71 21.682 249.792 21.71 ;
      END
   END FE_OFN6610_n_140234

   PIN FE_OFN6660_n_41611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.066 249.792 14.094 ;
      END
   END FE_OFN6660_n_41611

   PIN FE_OFN6723_n_41706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 179.698 0.0 179.726 0.163 ;
      END
   END FE_OFN6723_n_41706

   PIN FE_OFN6734_n_41994
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.474 249.792 55.502 ;
      END
   END FE_OFN6734_n_41994

   PIN FE_OFN6770_n_143423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.946 0.0 224.974 0.163 ;
      END
   END FE_OFN6770_n_143423

   PIN FE_OFN6842_n_41015
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.33 249.792 41.358 ;
      END
   END FE_OFN6842_n_41015

   PIN FE_OFN6876_n_41734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 41.202 249.792 41.23 ;
      END
   END FE_OFN6876_n_41734

   PIN FE_OFN6961_n_140210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.41 249.792 55.438 ;
      END
   END FE_OFN6961_n_140210

   PIN FE_OFN7004_n_140202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.85 0.0 204.878 0.163 ;
      END
   END FE_OFN7004_n_140202

   PIN FE_OFN7022_n_66979
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 230.514 0.0 230.542 0.163 ;
      END
   END FE_OFN7022_n_66979

   PIN FE_OFN8169_n_26637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.45 117.597 230.478 117.76 ;
      END
   END FE_OFN8169_n_26637

   PIN FE_OFN8329_n_31307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.362 0.0 181.39 0.163 ;
      END
   END FE_OFN8329_n_31307

   PIN FE_OFN8463_n_25371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.962 249.792 62.99 ;
      END
   END FE_OFN8463_n_25371

   PIN FE_OFN8477_n_30279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.386 0.0 230.414 0.163 ;
      END
   END FE_OFN8477_n_30279

   PIN FE_OFN8491_n_29557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.25 0.0 211.278 0.163 ;
      END
   END FE_OFN8491_n_29557

   PIN FE_OFN8577_n_29968
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.81 0.0 245.838 0.163 ;
      END
   END FE_OFN8577_n_29968

   PIN FE_OFN8703_n_31118
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 19.314 249.792 19.342 ;
      END
   END FE_OFN8703_n_31118

   PIN FE_OFN8799_n_25382
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.986 0.0 192.014 0.163 ;
      END
   END FE_OFN8799_n_25382

   PIN FE_OFN9238_delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.362 0.0 197.39 0.163 ;
      END
   END FE_OFN9238_delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_

   PIN FE_OFN9464_b_7_8_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.226 249.792 26.254 ;
      END
   END FE_OFN9464_b_7_8_11

   PIN FE_OFN9467_b_7_8_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.762 249.792 11.79 ;
      END
   END FE_OFN9467_b_7_8_10

   PIN FE_OFN9480_b_7_8_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.362 249.792 21.39 ;
      END
   END FE_OFN9480_b_7_8_5

   PIN FE_OFN9486_b_7_8_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 25.842 249.792 25.87 ;
      END
   END FE_OFN9486_b_7_8_3

   PIN FE_OFN9489_b_7_8_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.226 249.792 18.254 ;
      END
   END FE_OFN9489_b_7_8_2

   PIN FE_OFN9557_b_7_6_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.466 249.792 52.494 ;
      END
   END FE_OFN9557_b_7_6_6

   PIN FE_OFN9563_b_7_6_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 75.186 249.792 75.214 ;
      END
   END FE_OFN9563_b_7_6_5

   PIN FE_OFN9566_b_7_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 19.25 249.792 19.278 ;
      END
   END FE_OFN9566_b_7_6_4

   PIN FE_OFN9568_b_7_6_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.53 249.792 44.558 ;
      END
   END FE_OFN9568_b_7_6_3

   PIN FE_OFN9573_b_7_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 59.954 249.792 59.982 ;
      END
   END FE_OFN9573_b_7_6_2

   PIN FE_OFN9575_b_7_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.562 249.792 40.59 ;
      END
   END FE_OFN9575_b_7_6_2

   PIN FE_OFN9576_b_7_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.274 117.597 220.302 117.76 ;
      END
   END FE_OFN9576_b_7_6_1

   PIN FE_OFN9580_b_7_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 19.122 249.792 19.15 ;
      END
   END FE_OFN9580_b_7_6_0

   PIN FE_OFN9732_b_7_0_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.282 249.792 55.31 ;
      END
   END FE_OFN9732_b_7_0_10

   PIN FE_OFN9735_b_7_0_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 55.666 249.792 55.694 ;
      END
   END FE_OFN9735_b_7_0_9

   PIN FE_OFN9752_b_7_0_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 60.274 249.792 60.302 ;
      END
   END FE_OFN9752_b_7_0_5

   PIN FE_OFN9757_b_7_0_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.986 249.792 56.014 ;
      END
   END FE_OFN9757_b_7_0_4

   PIN FE_OFN9765_b_7_0_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 62.45 249.792 62.478 ;
      END
   END FE_OFN9765_b_7_0_2

   PIN FE_OFN9769_b_7_0_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.754 249.792 40.782 ;
      END
   END FE_OFN9769_b_7_0_1

   PIN FE_OFN9772_b_7_0_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.682 249.792 29.71 ;
      END
   END FE_OFN9772_b_7_0_0

   PIN FE_OFN9858_b_4_8_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.17 0.0 61.198 0.163 ;
      END
   END FE_OFN9858_b_4_8_13

   PIN FE_OFN9860_b_4_8_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 68.018 0.0 68.046 0.163 ;
      END
   END FE_OFN9860_b_4_8_12

   PIN FE_OFN9862_b_4_8_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.17 0.0 69.198 0.163 ;
      END
   END FE_OFN9862_b_4_8_11

   PIN FE_OFN9883_b_4_8_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.258 0.0 78.286 0.082 ;
      END
   END FE_OFN9883_b_4_8_2

   PIN FE_OFN9961_b_4_6_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.026 0.0 79.054 0.082 ;
      END
   END FE_OFN9961_b_4_6_3

   PIN FE_OFN9964_b_4_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.058 0.0 83.086 0.082 ;
      END
   END FE_OFN9964_b_4_6_2

   PIN b_4_8_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.858 117.597 103.886 117.76 ;
      END
   END b_4_8_3

   PIN b_7_0_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.322 249.792 70.35 ;
      END
   END b_7_0_7

   PIN b_7_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 56.05 249.792 56.078 ;
      END
   END b_7_6_0

   PIN b_7_6_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.146 117.597 204.174 117.76 ;
      END
   END b_7_6_10

   PIN b_7_6_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 218.802 117.597 218.83 117.76 ;
      END
   END b_7_6_11

   PIN b_7_6_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 222.834 117.597 222.862 117.76 ;
      END
   END b_7_6_14

   PIN b_7_6_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 215.218 117.597 215.246 117.76 ;
      END
   END b_7_6_15

   PIN b_7_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.546 117.597 226.574 117.76 ;
      END
   END b_7_6_4

   PIN b_7_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.578 249.792 62.606 ;
      END
   END b_7_6_7

   PIN b_7_6_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 218.994 117.597 219.022 117.76 ;
      END
   END b_7_6_9

   PIN b_7_8_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 170.482 117.597 170.51 117.76 ;
      END
   END b_7_8_7

   PIN b_7_8_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 196.146 117.597 196.174 117.76 ;
      END
   END b_7_8_8

   PIN delay_mul_ln34_unr7_unr8_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 174.578 0.0 174.606 0.163 ;
      END
   END delay_mul_ln34_unr7_unr8_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.114 0.0 96.142 0.163 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr8_unr7_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 173.234 0.0 173.262 0.163 ;
      END
   END delay_mul_ln34_unr8_unr7_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr8_unr7_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.458 0.0 169.486 0.163 ;
      END
   END delay_mul_ln34_unr8_unr7_stage2_stallmux_z_3_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 243.314 117.597 243.342 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.066 117.597 246.094 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.002 117.597 246.03 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_3_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.57 117.678 107.598 117.76 ;
      END
   END ispd_clk

   PIN mul_4647_72_n_181
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.322 0.163 62.35 ;
      END
   END mul_4647_72_n_181

   PIN mul_4647_72_n_182
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.282 0.0 15.31 0.163 ;
      END
   END mul_4647_72_n_182

   PIN mul_4647_72_n_53
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.562 0.163 40.59 ;
      END
   END mul_4647_72_n_53

   PIN mul_4647_72_n_69
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.33 0.163 33.358 ;
      END
   END mul_4647_72_n_69

   PIN mul_4647_72_n_779
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.266 0.163 33.294 ;
      END
   END mul_4647_72_n_779

   PIN mul_4649_72_n_825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.458 0.0 121.486 0.163 ;
      END
   END mul_4649_72_n_825

   PIN mul_4649_72_n_88
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.25 0.0 115.278 0.163 ;
      END
   END mul_4649_72_n_88

   PIN mul_4651_72_n_285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.322 0.0 94.35 0.163 ;
      END
   END mul_4651_72_n_285

   PIN mul_4664_72_n_241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.674 0.0 74.702 0.163 ;
      END
   END mul_4664_72_n_241

   PIN mul_4664_72_n_242
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.762 0.0 75.79 0.163 ;
      END
   END mul_4664_72_n_242

   PIN mul_4664_72_n_317
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.754 0.0 56.782 0.163 ;
      END
   END mul_4664_72_n_317

   PIN mul_4664_72_n_318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.69 0.0 56.718 0.163 ;
      END
   END mul_4664_72_n_318

   PIN mul_4664_72_n_319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.642 0.0 54.67 0.163 ;
      END
   END mul_4664_72_n_319

   PIN mul_4664_72_n_813
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.202 0.0 33.23 0.163 ;
      END
   END mul_4664_72_n_813

   PIN mul_4664_72_n_825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.322 0.0 62.35 0.163 ;
      END
   END mul_4664_72_n_825

   PIN mul_4664_72_n_84
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.202 0.0 65.23 0.163 ;
      END
   END mul_4664_72_n_84

   PIN mul_4664_72_n_848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.498 0.0 32.526 0.163 ;
      END
   END mul_4664_72_n_848

   PIN mul_4664_72_n_85
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.41 0.0 71.438 0.163 ;
      END
   END mul_4664_72_n_85

   PIN mul_4664_72_n_88
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.746 0.0 37.774 0.163 ;
      END
   END mul_4664_72_n_88

   PIN mul_4698_72_n_100
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.954 249.792 3.982 ;
      END
   END mul_4698_72_n_100

   PIN mul_4698_72_n_99
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.698 249.792 3.726 ;
      END
   END mul_4698_72_n_99

   PIN mul_4700_72_n_178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.706 249.792 6.734 ;
      END
   END mul_4700_72_n_178

   PIN mul_4700_72_n_179
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.634 249.792 3.662 ;
      END
   END mul_4700_72_n_179

   PIN n_101492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 161.458 0.0 161.486 0.163 ;
      END
   END n_101492

   PIN n_102695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.77 249.792 110.798 ;
      END
   END n_102695

   PIN n_103071
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.026 117.597 215.054 117.76 ;
      END
   END n_103071

   PIN n_103939
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 225.458 117.597 225.486 117.76 ;
      END
   END n_103939

   PIN n_103940
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.218 117.597 215.246 117.76 ;
      END
   END n_103940

   PIN n_106720
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.706 249.792 110.734 ;
      END
   END n_106720

   PIN n_107989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.946 0.0 40.974 0.163 ;
      END
   END n_107989

   PIN n_108267
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.634 117.597 203.662 117.76 ;
      END
   END n_108267

   PIN n_108268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.41 117.597 207.438 117.76 ;
      END
   END n_108268

   PIN n_108688
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.018 117.597 196.046 117.76 ;
      END
   END n_108688

   PIN n_110443
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 60.21 249.792 60.238 ;
      END
   END n_110443

   PIN n_110533
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 90.482 249.792 90.51 ;
      END
   END n_110533

   PIN n_112122
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.202 0.163 33.23 ;
      END
   END n_112122

   PIN n_112183
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.482 0.0 66.51 0.082 ;
      END
   END n_112183

   PIN n_112413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.138 0.0 97.166 0.163 ;
      END
   END n_112413

   PIN n_112659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.866 0.0 74.894 0.163 ;
      END
   END n_112659

   PIN n_114178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.714 0.0 49.742 0.163 ;
      END
   END n_114178

   PIN n_114182
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.594 0.0 12.622 0.163 ;
      END
   END n_114182

   PIN n_114494
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.738 0.0 26.766 0.163 ;
      END
   END n_114494

   PIN n_114496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.674 0.0 26.702 0.163 ;
      END
   END n_114496

   PIN n_114524
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.658 0.0 12.686 0.163 ;
      END
   END n_114524

   PIN n_114615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.546 0.0 42.574 0.163 ;
      END
   END n_114615

   PIN n_114617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.058 0.0 19.086 0.163 ;
      END
   END n_114617

   PIN n_114672
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.69 117.597 48.718 117.76 ;
      END
   END n_114672

   PIN n_114673
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.866 0.0 26.894 0.163 ;
      END
   END n_114673

   PIN n_114676
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.058 0.0 19.086 0.163 ;
      END
   END n_114676

   PIN n_114855
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.89 0.0 43.918 0.163 ;
      END
   END n_114855

   PIN n_114920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.866 0.0 58.894 0.163 ;
      END
   END n_114920

   PIN n_114921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.674 0.0 58.702 0.163 ;
      END
   END n_114921

   PIN n_115152
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.402 0.0 52.43 0.163 ;
      END
   END n_115152

   PIN n_115153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.21 0.0 52.238 0.163 ;
      END
   END n_115153

   PIN n_115190
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.594 0.0 44.622 0.163 ;
      END
   END n_115190

   PIN n_115308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.554 0.0 13.582 0.163 ;
      END
   END n_115308

   PIN n_115309
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.754 0.0 16.782 0.163 ;
      END
   END n_115309

   PIN n_115311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.418 0.0 50.446 0.163 ;
      END
   END n_115311

   PIN n_115543
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.994 0.0 19.022 0.163 ;
      END
   END n_115543

   PIN n_115582
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.642 0.0 30.67 0.163 ;
      END
   END n_115582

   PIN n_115593
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.786 0.0 20.814 0.163 ;
      END
   END n_115593

   PIN n_115606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.754 0.0 48.782 0.163 ;
      END
   END n_115606

   PIN n_115661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.034 0.0 50.062 0.163 ;
      END
   END n_115661

   PIN n_115793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.938 0.0 45.966 0.163 ;
      END
   END n_115793

   PIN n_115794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 46.13 0.0 46.158 0.163 ;
      END
   END n_115794

   PIN n_115810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.57 0.0 11.598 0.163 ;
      END
   END n_115810

   PIN n_116281
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.802 0.0 26.83 0.163 ;
      END
   END n_116281

   PIN n_116796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.802 0.0 34.83 0.163 ;
      END
   END n_116796

   PIN n_117132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.722 0.0 76.75 0.163 ;
      END
   END n_117132

   PIN n_117734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.122 0.0 19.15 0.163 ;
      END
   END n_117734

   PIN n_117835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.418 0.0 34.446 0.163 ;
      END
   END n_117835

   PIN n_118212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.346 0.0 47.374 0.163 ;
      END
   END n_118212

   PIN n_118398
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.306 0.0 16.334 0.163 ;
      END
   END n_118398

   PIN n_119074
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.162 0.163 114.19 ;
      END
   END n_119074

   PIN n_120882
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.538 117.597 47.566 117.76 ;
      END
   END n_120882

   PIN n_121314
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.866 0.0 26.894 0.163 ;
      END
   END n_121314

   PIN n_121751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.706 0.0 30.734 0.163 ;
      END
   END n_121751

   PIN n_121989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.034 0.0 26.062 0.163 ;
      END
   END n_121989

   PIN n_122315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.706 0.0 22.734 0.163 ;
      END
   END n_122315

   PIN n_122349
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.578 0.0 30.606 0.163 ;
      END
   END n_122349

   PIN n_123446
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.034 0.0 42.062 0.163 ;
      END
   END n_123446

   PIN n_124498
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.602 0.163 47.63 ;
      END
   END n_124498

   PIN n_124539
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.682 117.597 37.71 117.76 ;
      END
   END n_124539

   PIN n_124540
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.946 117.597 40.974 117.76 ;
      END
   END n_124540

   PIN n_124638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.562 0.0 16.59 0.163 ;
      END
   END n_124638

   PIN n_124639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.986 0.0 24.014 0.163 ;
      END
   END n_124639

   PIN n_125192
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.666 0.163 71.694 ;
      END
   END n_125192

   PIN n_125461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.026 0.0 23.054 0.163 ;
      END
   END n_125461

   PIN n_125695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.466 0.163 52.494 ;
      END
   END n_125695

   PIN n_125716
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.49 0.0 13.518 0.163 ;
      END
   END n_125716

   PIN n_127036
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.498 0.0 16.526 0.163 ;
      END
   END n_127036

   PIN n_127040
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.93 0.0 26.958 0.163 ;
      END
   END n_127040

   PIN n_127190
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.922 117.597 47.95 117.76 ;
      END
   END n_127190

   PIN n_127195
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.682 0.0 13.71 0.163 ;
      END
   END n_127195

   PIN n_127589
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.402 0.163 52.43 ;
      END
   END n_127589

   PIN n_127666
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.866 0.163 90.894 ;
      END
   END n_127666

   PIN n_128129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.274 0.0 28.302 0.163 ;
      END
   END n_128129

   PIN n_128287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.786 0.163 44.814 ;
      END
   END n_128287

   PIN n_128296
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.794 0.0 7.822 0.163 ;
      END
   END n_128296

   PIN n_128768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.01 117.597 57.038 117.76 ;
      END
   END n_128768

   PIN n_129724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.722 0.163 44.75 ;
      END
   END n_129724

   PIN n_130012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.77 0.0 22.798 0.163 ;
      END
   END n_130012

   PIN n_130016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.434 0.0 16.462 0.163 ;
      END
   END n_130016

   PIN n_131230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.882 0.0 24.91 0.163 ;
      END
   END n_131230

   PIN n_132777
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.93 117.597 26.958 117.76 ;
      END
   END n_132777

   PIN n_133344
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.818 0.0 16.846 0.163 ;
      END
   END n_133344

   PIN n_133767
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.45 0.0 38.478 0.163 ;
      END
   END n_133767

   PIN n_137225
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.874 0.0 45.902 0.163 ;
      END
   END n_137225

   PIN n_137233
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.186 249.792 11.214 ;
      END
   END n_137233

   PIN n_137728
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.682 0.0 181.71 0.163 ;
      END
   END n_137728

   PIN n_137826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 87.218 249.792 87.246 ;
      END
   END n_137826

   PIN n_137827
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.634 0.0 107.662 0.163 ;
      END
   END n_137827

   PIN n_137828
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.586 0.0 57.614 0.163 ;
      END
   END n_137828

   PIN n_137851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.098 0.0 42.126 0.163 ;
      END
   END n_137851

   PIN n_140213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 232.626 0.0 232.654 0.163 ;
      END
   END n_140213

   PIN n_142851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.618 0.0 61.646 0.082 ;
      END
   END n_142851

   PIN n_142964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.266 0.0 65.294 0.163 ;
      END
   END n_142964

   PIN n_143483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 234.418 0.0 234.446 0.082 ;
      END
   END n_143483

   PIN n_143496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 17.522 249.792 17.55 ;
      END
   END n_143496

   PIN n_143630
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.714 249.792 33.742 ;
      END
   END n_143630

   PIN n_143743
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.562 0.163 48.59 ;
      END
   END n_143743

   PIN n_143933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.57 0.0 107.598 0.163 ;
      END
   END n_143933

   PIN n_144109
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 84.53 0.0 84.558 0.163 ;
      END
   END n_144109

   PIN n_144135
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.802 117.597 218.83 117.76 ;
      END
   END n_144135

   PIN n_144158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.978 249.792 45.006 ;
      END
   END n_144158

   PIN n_24056
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.794 0.0 199.822 0.163 ;
      END
   END n_24056

   PIN n_25134
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.01 0.0 169.038 0.163 ;
      END
   END n_25134

   PIN n_25376
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.69 249.792 40.718 ;
      END
   END n_25376

   PIN n_26011
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.506 0.0 203.534 0.163 ;
      END
   END n_26011

   PIN n_26383
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.13 117.597 150.158 117.76 ;
      END
   END n_26383

   PIN n_26633
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 60.146 249.792 60.174 ;
      END
   END n_26633

   PIN n_27338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.618 117.597 109.646 117.76 ;
      END
   END n_27338

   PIN n_27740
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.93 117.597 106.958 117.76 ;
      END
   END n_27740

   PIN n_27741
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.802 117.597 106.83 117.76 ;
      END
   END n_27741

   PIN n_28380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.09 0.0 215.118 0.163 ;
      END
   END n_28380

   PIN n_28496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.834 249.792 94.862 ;
      END
   END n_28496

   PIN n_28631
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.354 0.0 42.382 0.163 ;
      END
   END n_28631

   PIN n_28640
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.354 0.0 186.382 0.163 ;
      END
   END n_28640

   PIN n_28780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 99.058 249.792 99.086 ;
      END
   END n_28780

   PIN n_29125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 213.042 0.0 213.07 0.163 ;
      END
   END n_29125

   PIN n_31876
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.602 0.0 103.63 0.163 ;
      END
   END n_31876

   PIN n_33226
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.09 0.0 47.118 0.163 ;
      END
   END n_33226

   PIN n_33292
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.074 0.0 97.102 0.163 ;
      END
   END n_33292

   PIN n_33293
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.338 0.0 84.366 0.163 ;
      END
   END n_33293

   PIN n_33375
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.514 0.0 62.542 0.163 ;
      END
   END n_33375

   PIN n_33782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.466 0.0 84.494 0.163 ;
      END
   END n_33782

   PIN n_34260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 238.13 0.0 238.158 0.163 ;
      END
   END n_34260

   PIN n_34345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.97 0.0 73.998 0.163 ;
      END
   END n_34345

   PIN n_35072
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.49 0.0 69.518 0.163 ;
      END
   END n_35072

   PIN n_35096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.722 0.0 116.75 0.163 ;
      END
   END n_35096

   PIN n_36000
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.394 0.0 73.422 0.163 ;
      END
   END n_36000

   PIN n_36612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.122 0.0 75.15 0.163 ;
      END
   END n_36612

   PIN n_37235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.122 0.0 59.15 0.163 ;
      END
   END n_37235

   PIN n_37476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.954 0.0 67.982 0.163 ;
      END
   END n_37476

   PIN n_40827
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.226 0.0 162.254 0.163 ;
      END
   END n_40827

   PIN n_40897
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 232.498 0.0 232.526 0.163 ;
      END
   END n_40897

   PIN n_40960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.578 249.792 6.606 ;
      END
   END n_40960

   PIN n_41417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 2.482 249.792 2.51 ;
      END
   END n_41417

   PIN n_41500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.57 249.792 3.598 ;
      END
   END n_41500

   PIN n_41612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.994 249.792 19.022 ;
      END
   END n_41612

   PIN n_41734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.618 249.792 29.646 ;
      END
   END n_41734

   PIN n_41834
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.506 249.792 3.534 ;
      END
   END n_41834

   PIN n_41962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 13.874 249.792 13.902 ;
      END
   END n_41962

   PIN n_42268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.938 249.792 77.966 ;
      END
   END n_42268

   PIN n_42269
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.874 249.792 77.902 ;
      END
   END n_42269

   PIN n_42354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 98.482 249.792 98.51 ;
      END
   END n_42354

   PIN n_42362
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 105.97 249.792 105.998 ;
      END
   END n_42362

   PIN n_42412
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.81 249.792 77.838 ;
      END
   END n_42412

   PIN n_42413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.746 249.792 77.774 ;
      END
   END n_42413

   PIN n_42443
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.866 249.792 106.894 ;
      END
   END n_42443

   PIN n_42504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 79.09 249.792 79.118 ;
      END
   END n_42504

   PIN n_42506
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 98.226 249.792 98.254 ;
      END
   END n_42506

   PIN n_42608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.642 249.792 102.67 ;
      END
   END n_42608

   PIN n_42807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.45 249.792 110.478 ;
      END
   END n_42807

   PIN n_42921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.514 249.792 94.542 ;
      END
   END n_42921

   PIN n_43096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.514 249.792 14.542 ;
      END
   END n_43096

   PIN n_43134
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.89 249.792 99.918 ;
      END
   END n_43134

   PIN n_43240
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.506 249.792 99.534 ;
      END
   END n_43240

   PIN n_43320
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.922 249.792 55.95 ;
      END
   END n_43320

   PIN n_43384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 114.162 249.792 114.19 ;
      END
   END n_43384

   PIN n_43416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.45 249.792 94.478 ;
      END
   END n_43416

   PIN n_43545
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 68.018 249.792 68.046 ;
      END
   END n_43545

   PIN n_43643
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.386 249.792 94.414 ;
      END
   END n_43643

   PIN n_43707
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.13 249.792 110.158 ;
      END
   END n_43707

   PIN n_44058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 98.098 249.792 98.126 ;
      END
   END n_44058

   PIN n_44137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.674 117.597 226.702 117.76 ;
      END
   END n_44137

   PIN n_44356
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.93 249.792 18.958 ;
      END
   END n_44356

   PIN n_44415
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.258 249.792 70.286 ;
      END
   END n_44415

   PIN n_44594
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.826 249.792 99.854 ;
      END
   END n_44594

   PIN n_44658
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.442 249.792 99.47 ;
      END
   END n_44658

   PIN n_45114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 105.906 249.792 105.934 ;
      END
   END n_45114

   PIN n_45130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.194 249.792 70.222 ;
      END
   END n_45130

   PIN n_45297
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 67.698 249.792 67.726 ;
      END
   END n_45297

   PIN n_45432
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.162 249.792 26.19 ;
      END
   END n_45432

   PIN n_45433
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.098 249.792 26.126 ;
      END
   END n_45433

   PIN n_45435
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.786 249.792 52.814 ;
      END
   END n_45435

   PIN n_45598
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 91.762 249.792 91.79 ;
      END
   END n_45598

   PIN n_45795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.85 249.792 84.878 ;
      END
   END n_45795

   PIN n_45796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 84.722 249.792 84.75 ;
      END
   END n_45796

   PIN n_46004
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 28.914 249.792 28.942 ;
      END
   END n_46004

   PIN n_46071
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.554 249.792 29.582 ;
      END
   END n_46071

   PIN n_46080
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.362 249.792 37.39 ;
      END
   END n_46080

   PIN n_46178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.322 0.0 86.35 0.163 ;
      END
   END n_46178

   PIN n_46181
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.002 249.792 30.03 ;
      END
   END n_46181

   PIN n_46217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 67.634 249.792 67.662 ;
      END
   END n_46217

   PIN n_46227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.298 249.792 37.326 ;
      END
   END n_46227

   PIN n_46333
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.242 249.792 48.27 ;
      END
   END n_46333

   PIN n_46334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.514 249.792 6.542 ;
      END
   END n_46334

   PIN n_46340
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 25.97 249.792 25.998 ;
      END
   END n_46340

   PIN n_46341
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 25.906 249.792 25.934 ;
      END
   END n_46341

   PIN n_46365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.45 249.792 6.478 ;
      END
   END n_46365

   PIN n_46513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.49 249.792 29.518 ;
      END
   END n_46513

   PIN n_46588
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.522 249.792 33.55 ;
      END
   END n_46588

   PIN n_46658
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.698 249.792 11.726 ;
      END
   END n_46658

   PIN n_46660
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 17.778 249.792 17.806 ;
      END
   END n_46660

   PIN n_46774
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.386 249.792 6.414 ;
      END
   END n_46774

   PIN n_46851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 67.954 249.792 67.982 ;
      END
   END n_46851

   PIN n_46932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.65 249.792 33.678 ;
      END
   END n_46932

   PIN n_46954
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 47.666 249.792 47.694 ;
      END
   END n_46954

   PIN n_47028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.474 0.0 247.502 0.163 ;
      END
   END n_47028

   PIN n_47607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.386 0.0 62.414 0.163 ;
      END
   END n_47607

   PIN n_47644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.442 249.792 3.47 ;
      END
   END n_47644

   PIN n_47750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.826 0.0 83.854 0.163 ;
      END
   END n_47750

   PIN n_47929
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.714 0.0 57.742 0.163 ;
      END
   END n_47929

   PIN n_48546
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.618 249.792 37.646 ;
      END
   END n_48546

   PIN n_48611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.85 0.0 44.878 0.163 ;
      END
   END n_48611

   PIN n_48880
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.554 249.792 37.582 ;
      END
   END n_48880

   PIN n_48997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.426 249.792 29.454 ;
      END
   END n_48997

   PIN n_49055
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.362 249.792 29.39 ;
      END
   END n_49055

   PIN n_49568
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.794 0.0 7.822 0.163 ;
      END
   END n_49568

   PIN n_49769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 3.442 249.792 3.47 ;
      END
   END n_49769

   PIN n_49987
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.13 249.792 70.158 ;
      END
   END n_49987

   PIN n_50107
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.322 249.792 6.35 ;
      END
   END n_50107

   PIN n_50238
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.322 249.792 102.35 ;
      END
   END n_50238

   PIN n_50246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 79.41 249.792 79.438 ;
      END
   END n_50246

   PIN n_50397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 17.65 249.792 17.678 ;
      END
   END n_50397

   PIN n_50495
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.386 249.792 110.414 ;
      END
   END n_50495

   PIN n_50522
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.634 249.792 99.662 ;
      END
   END n_50522

   PIN n_50818
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 91.954 249.792 91.982 ;
      END
   END n_50818

   PIN n_50937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.666 0.0 191.694 0.163 ;
      END
   END n_50937

   PIN n_51078
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 67.57 249.792 67.598 ;
      END
   END n_51078

   PIN n_51110
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.034 249.792 26.062 ;
      END
   END n_51110

   PIN n_51111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 25.842 249.792 25.87 ;
      END
   END n_51111

   PIN n_51211
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.01 249.792 33.038 ;
      END
   END n_51211

   PIN n_51212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.946 249.792 32.974 ;
      END
   END n_51212

   PIN n_51988
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 67.89 249.792 67.918 ;
      END
   END n_51988

   PIN n_52066
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.602 0.0 191.63 0.163 ;
      END
   END n_52066

   PIN n_52279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 79.282 249.792 79.31 ;
      END
   END n_52279

   PIN n_52455
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.106 249.792 77.134 ;
      END
   END n_52455

   PIN n_52456
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 76.978 249.792 77.006 ;
      END
   END n_52456

   PIN n_52502
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 33.33 249.792 33.358 ;
      END
   END n_52502

   PIN n_52697
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.066 249.792 110.094 ;
      END
   END n_52697

   PIN n_52749
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.258 249.792 102.286 ;
      END
   END n_52749

   PIN n_52750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.802 249.792 106.83 ;
      END
   END n_52750

   PIN n_52873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 98.162 249.792 98.19 ;
      END
   END n_52873

   PIN n_52994
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.346 249.792 55.374 ;
      END
   END n_52994

   PIN n_53090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 2.802 249.792 2.83 ;
      END
   END n_53090

   PIN n_53725
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.514 249.792 102.542 ;
      END
   END n_53725

   PIN n_53750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.57 249.792 99.598 ;
      END
   END n_53750

   PIN n_53835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.786 0.0 44.814 0.163 ;
      END
   END n_53835

   PIN n_54049
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.298 249.792 29.326 ;
      END
   END n_54049

   PIN n_54060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 15.41 249.792 15.438 ;
      END
   END n_54060

   PIN n_54354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 13.81 249.792 13.838 ;
      END
   END n_54354

   PIN n_54357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.634 249.792 11.662 ;
      END
   END n_54357

   PIN n_54358
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 11.122 249.792 11.15 ;
      END
   END n_54358

   PIN n_54853
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 190.578 0.0 190.606 0.163 ;
      END
   END n_54853

   PIN n_54873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 113.842 249.792 113.87 ;
      END
   END n_54873

   PIN n_54905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.194 249.792 110.222 ;
      END
   END n_54905

   PIN n_54906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.098 117.597 242.126 117.76 ;
      END
   END n_54906

   PIN n_54932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 234.354 117.597 234.382 117.76 ;
      END
   END n_54932

   PIN n_54940
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.674 249.792 106.702 ;
      END
   END n_54940

   PIN n_54943
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.61 117.597 226.638 117.76 ;
      END
   END n_54943

   PIN n_54953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.762 249.792 99.79 ;
      END
   END n_54953

   PIN n_55031
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.914 249.792 44.942 ;
      END
   END n_55031

   PIN n_55096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.81 249.792 21.838 ;
      END
   END n_55096

   PIN n_55097
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.746 249.792 21.774 ;
      END
   END n_55097

   PIN n_5512
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.378 0.0 19.406 0.163 ;
      END
   END n_5512

   PIN n_55141
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.938 117.597 245.966 117.76 ;
      END
   END n_55141

   PIN n_55158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.49 249.792 37.518 ;
      END
   END n_55158

   PIN n_55332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 91.89 249.792 91.918 ;
      END
   END n_55332

   PIN n_55444
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.682 249.792 21.71 ;
      END
   END n_55444

   PIN n_55445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 21.81 249.792 21.838 ;
      END
   END n_55445

   PIN n_55540
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 157.554 0.0 157.582 0.163 ;
      END
   END n_55540

   PIN n_55560
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 78.962 249.792 78.99 ;
      END
   END n_55560

   PIN n_55599
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.882 249.792 32.91 ;
      END
   END n_55599

   PIN n_55648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.994 0.0 147.022 0.163 ;
      END
   END n_55648

   PIN n_55722
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.146 0.0 140.174 0.163 ;
      END
   END n_55722

   PIN n_55790
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 9.778 249.792 9.806 ;
      END
   END n_55790

   PIN n_5584
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.802 0.0 10.83 0.163 ;
      END
   END n_5584

   PIN n_55908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.042 249.792 45.07 ;
      END
   END n_55908

   PIN n_56447
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.322 249.792 110.35 ;
      END
   END n_56447

   PIN n_56448
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.258 249.792 110.286 ;
      END
   END n_56448

   PIN n_56512
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 40.818 249.792 40.846 ;
      END
   END n_56512

   PIN n_56516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.074 249.792 41.102 ;
      END
   END n_56516

   PIN n_56956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 187.762 0.0 187.79 0.163 ;
      END
   END n_56956

   PIN n_57348
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 33.266 249.792 33.294 ;
      END
   END n_57348

   PIN n_57368
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 56.242 249.792 56.27 ;
      END
   END n_57368

   PIN n_57417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.138 249.792 33.166 ;
      END
   END n_57417

   PIN n_57444
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.73 0.0 199.758 0.163 ;
      END
   END n_57444

   PIN n_57615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.338 249.792 92.366 ;
      END
   END n_57615

   PIN n_57620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.394 0.0 65.422 0.163 ;
      END
   END n_57620

   PIN n_57624
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.938 249.792 29.966 ;
      END
   END n_57624

   PIN n_57629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.946 249.792 40.974 ;
      END
   END n_57629

   PIN n_57726
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.874 0.0 245.902 0.163 ;
      END
   END n_57726

   PIN n_57746
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 36.786 249.792 36.814 ;
      END
   END n_57746

   PIN n_57903
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.138 117.597 113.166 117.76 ;
      END
   END n_57903

   PIN n_57935
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.234 249.792 37.262 ;
      END
   END n_57935

   PIN n_57983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.21 117.597 164.238 117.76 ;
      END
   END n_57983

   PIN n_58082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 106.546 249.792 106.574 ;
      END
   END n_58082

   PIN n_58177
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 110.002 249.792 110.03 ;
      END
   END n_58177

   PIN n_58261
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 222.77 117.597 222.798 117.76 ;
      END
   END n_58261

   PIN n_58290
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.402 117.597 220.43 117.76 ;
      END
   END n_58290

   PIN n_58294
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.338 117.597 220.366 117.76 ;
      END
   END n_58294

   PIN n_58385
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 21.554 249.792 21.582 ;
      END
   END n_58385

   PIN n_58399
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.49 249.792 21.518 ;
      END
   END n_58399

   PIN n_58400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 21.426 249.792 21.454 ;
      END
   END n_58400

   PIN n_58672
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 242.034 0.0 242.062 0.163 ;
      END
   END n_58672

   PIN n_58674
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 13.746 249.792 13.774 ;
      END
   END n_58674

   PIN n_59053
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.85 249.792 44.878 ;
      END
   END n_59053

   PIN n_59056
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.786 249.792 44.814 ;
      END
   END n_59056

   PIN n_59131
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 18.162 249.792 18.19 ;
      END
   END n_59131

   PIN n_59166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.874 117.597 245.902 117.76 ;
      END
   END n_59166

   PIN n_59286
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.194 117.597 238.222 117.76 ;
      END
   END n_59286

   PIN n_59394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.762 117.597 163.79 117.76 ;
      END
   END n_59394

   PIN n_59605
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.858 0.0 143.886 0.163 ;
      END
   END n_59605

   PIN n_60089
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.546 117.597 130.574 117.76 ;
      END
   END n_60089

   PIN n_60346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.122 249.792 11.15 ;
      END
   END n_60346

   PIN n_60369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.474 0.0 207.502 0.163 ;
      END
   END n_60369

   PIN n_60370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.426 0.0 205.454 0.163 ;
      END
   END n_60370

   PIN n_60378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.066 249.792 70.094 ;
      END
   END n_60378

   PIN n_60427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.322 249.792 14.35 ;
      END
   END n_60427

   PIN n_60554
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 36.722 249.792 36.75 ;
      END
   END n_60554

   PIN n_60615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.626 249.792 40.654 ;
      END
   END n_60615

   PIN n_60632
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.466 249.792 44.494 ;
      END
   END n_60632

   PIN n_61085
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 29.234 249.792 29.262 ;
      END
   END n_61085

   PIN n_61149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.866 249.792 18.894 ;
      END
   END n_61149

   PIN n_61187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.002 249.792 14.03 ;
      END
   END n_61187

   PIN n_61461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.034 117.597 242.062 117.76 ;
      END
   END n_61461

   PIN n_61579
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 13.874 249.792 13.902 ;
      END
   END n_61579

   PIN n_61580
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.802 249.792 18.83 ;
      END
   END n_61580

   PIN n_61592
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.274 249.792 92.302 ;
      END
   END n_61592

   PIN n_61601
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.602 249.792 47.63 ;
      END
   END n_61601

   PIN n_61705
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.282 117.597 95.31 117.76 ;
      END
   END n_61705

   PIN n_61723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.522 0.0 57.55 0.163 ;
      END
   END n_61723

   PIN n_61755
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.834 0.0 102.862 0.163 ;
      END
   END n_61755

   PIN n_61873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.578 249.792 102.606 ;
      END
   END n_61873

   PIN n_61878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.13 117.597 238.158 117.76 ;
      END
   END n_61878

   PIN n_61893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.866 117.597 218.894 117.76 ;
      END
   END n_61893

   PIN n_61956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 9.714 249.792 9.742 ;
      END
   END n_61956

   PIN n_62290
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 13.618 249.792 13.646 ;
      END
   END n_62290

   PIN n_62406
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.458 249.792 41.486 ;
      END
   END n_62406

   PIN n_62437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.69 117.597 160.718 117.76 ;
      END
   END n_62437

   PIN n_62460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.314 117.597 211.342 117.76 ;
      END
   END n_62460

   PIN n_62694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 247.282 117.597 247.31 117.76 ;
      END
   END n_62694

   PIN n_62695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.514 117.597 230.542 117.76 ;
      END
   END n_62695

   PIN n_63124
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.162 249.792 18.19 ;
      END
   END n_63124

   PIN n_63132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.858 249.792 47.886 ;
      END
   END n_63132

   PIN n_63155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.394 0.0 89.422 0.163 ;
      END
   END n_63155

   PIN n_63260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 176.818 117.597 176.846 117.76 ;
      END
   END n_63260

   PIN n_63263
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 228.018 117.597 228.046 117.76 ;
      END
   END n_63263

   PIN n_63360
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.49 0.0 181.518 0.163 ;
      END
   END n_63360

   PIN n_63423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 21.874 249.792 21.902 ;
      END
   END n_63423

   PIN n_63445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.458 249.792 33.486 ;
      END
   END n_63445

   PIN n_63901
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.698 117.597 155.726 117.76 ;
      END
   END n_63901

   PIN n_64318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.042 117.597 149.07 117.76 ;
      END
   END n_64318

   PIN n_64366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.57 249.792 11.598 ;
      END
   END n_64366

   PIN n_64478
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 25.202 249.792 25.23 ;
      END
   END n_64478

   PIN n_64560
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.626 117.597 224.654 117.76 ;
      END
   END n_64560

   PIN n_64768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 9.842 249.792 9.87 ;
      END
   END n_64768

   PIN n_64772
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 44.722 249.792 44.75 ;
      END
   END n_64772

   PIN n_64912
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.938 117.597 149.966 117.76 ;
      END
   END n_64912

   PIN n_65026
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.562 117.597 224.59 117.76 ;
      END
   END n_65026

   PIN n_65319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.538 0.0 87.566 0.163 ;
      END
   END n_65319

   PIN n_65354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.962 117.597 142.99 117.76 ;
      END
   END n_65354

   PIN n_65426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.386 117.597 94.414 117.76 ;
      END
   END n_65426

   PIN n_65480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.794 249.792 47.822 ;
      END
   END n_65480

   PIN n_65483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.658 249.792 52.686 ;
      END
   END n_65483

   PIN n_65893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.402 249.792 52.43 ;
      END
   END n_65893

   PIN n_65894
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.338 249.792 52.366 ;
      END
   END n_65894

   PIN n_66724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 210.098 117.597 210.126 117.76 ;
      END
   END n_66724

   PIN n_66751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 52.274 249.792 52.302 ;
      END
   END n_66751

   PIN n_66842
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.786 249.792 84.814 ;
      END
   END n_66842

   PIN n_66843
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.722 249.792 84.75 ;
      END
   END n_66843

   PIN n_66867
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.978 117.597 149.006 117.76 ;
      END
   END n_66867

   PIN n_67068
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.17 0.0 125.198 0.163 ;
      END
   END n_67068

   PIN n_67215
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.73 249.792 47.758 ;
      END
   END n_67215

   PIN n_70345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.322 249.792 94.35 ;
      END
   END n_70345

   PIN n_70642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.706 249.792 94.734 ;
      END
   END n_70642

   PIN n_71222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.194 249.792 102.222 ;
      END
   END n_71222

   PIN n_71449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.442 0.0 99.47 0.163 ;
      END
   END n_71449

   PIN n_71795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.81 0.0 157.838 0.163 ;
      END
   END n_71795

   PIN n_77679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.45 0.0 134.478 0.163 ;
      END
   END n_77679

   PIN n_77842
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 46.194 0.0 46.222 0.163 ;
      END
   END n_77842

   PIN n_80858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.738 249.792 106.766 ;
      END
   END n_80858

   PIN n_81895
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.682 249.792 77.71 ;
      END
   END n_81895

   PIN n_82145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.594 117.597 180.622 117.76 ;
      END
   END n_82145

   PIN n_82355
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 79.026 249.792 79.054 ;
      END
   END n_82355

   PIN n_82437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 102.13 249.792 102.158 ;
      END
   END n_82437

   PIN n_8249
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.394 0.0 57.422 0.163 ;
      END
   END n_8249

   PIN n_82916
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.322 249.792 62.35 ;
      END
   END n_82916

   PIN n_83187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 91.826 249.792 91.854 ;
      END
   END n_83187

   PIN n_83203
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 79.346 249.792 79.374 ;
      END
   END n_83203

   PIN n_84332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 110.002 249.792 110.03 ;
      END
   END n_84332

   PIN n_85306
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 91.762 249.792 91.79 ;
      END
   END n_85306

   PIN n_85307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.77 249.792 94.798 ;
      END
   END n_85307

   PIN n_85541
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.402 0.0 180.43 0.163 ;
      END
   END n_85541

   PIN n_86195
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 59.826 249.792 59.854 ;
      END
   END n_86195

   PIN n_87554
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.69 117.597 176.718 117.76 ;
      END
   END n_87554

   PIN n_87555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.53 117.597 180.558 117.76 ;
      END
   END n_87555

   PIN n_88558
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 94.258 249.792 94.286 ;
      END
   END n_88558

   PIN n_95316
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 79.154 249.792 79.182 ;
      END
   END n_95316

   PIN n_95932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.162 0.0 42.19 0.163 ;
      END
   END n_95932

   PIN n_96299
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.034 117.597 186.062 117.76 ;
      END
   END n_96299

   PIN n_96642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.258 0.0 38.286 0.163 ;
      END
   END n_96642

   PIN n_97723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.682 0.0 149.71 0.163 ;
      END
   END n_97723

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER V1 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER M1 ;
         RECT 0.0 0.0 249.792 117.76 ;
   END
END h2_mgc_matrix_mult_a

MACRO h1_mgc_matrix_mult_a
   CLASS BLOCK ;
   FOREIGN h1 ;
   ORIGIN 0 0 ;
   SIZE 248.0 BY 154.88 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN15738_FE_OFN11549_n_142793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.714 154.717 113.742 154.88 ;
      END
   END FE_OCPN15738_FE_OFN11549_n_142793

   PIN FE_OFN10667_a_5_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 223.73 0.0 223.758 0.163 ;
      END
   END FE_OFN10667_a_5_6_4

   PIN FE_OFN10748_a_4_4_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 237.49 0.0 237.518 0.163 ;
      END
   END FE_OFN10748_a_4_4_4

   PIN FE_OFN10792_a_4_0_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.058 0.0 235.086 0.163 ;
      END
   END FE_OFN10792_a_4_0_5

   PIN FE_OFN10799_a_3_8_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 130.994 248.0 131.022 ;
      END
   END FE_OFN10799_a_3_8_7

   PIN FE_OFN10820_a_3_6_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 101.49 248.0 101.518 ;
      END
   END FE_OFN10820_a_3_6_7

   PIN FE_OFN10830_a_3_4_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.402 0.0 228.43 0.163 ;
      END
   END FE_OFN10830_a_3_4_5

   PIN FE_OFN10834_a_3_4_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 111.154 248.0 111.182 ;
      END
   END FE_OFN10834_a_3_4_0

   PIN FE_OFN10851_a_2_8_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 244.658 0.0 244.686 0.163 ;
      END
   END FE_OFN10851_a_2_8_4

   PIN FE_OFN10859_a_2_8_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 244.914 0.0 244.942 0.163 ;
      END
   END FE_OFN10859_a_2_8_1

   PIN FE_OFN10872_a_2_6_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 91.954 248.0 91.982 ;
      END
   END FE_OFN10872_a_2_6_7

   PIN FE_OFN10879_a_2_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.09 0.0 215.118 0.163 ;
      END
   END FE_OFN10879_a_2_6_4

   PIN FE_OFN10888_a_2_4_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 111.218 248.0 111.246 ;
      END
   END FE_OFN10888_a_2_4_7

   PIN FE_OFN10898_a_2_4_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.026 0.0 215.054 0.163 ;
      END
   END FE_OFN10898_a_2_4_1

   PIN FE_OFN10902_a_2_4_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 111.282 248.0 111.31 ;
      END
   END FE_OFN10902_a_2_4_0

   PIN FE_OFN10931_a_1_4_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 101.554 248.0 101.582 ;
      END
   END FE_OFN10931_a_1_4_0

   PIN FE_OFN10982_a_0_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 140.594 248.0 140.622 ;
      END
   END FE_OFN10982_a_0_6_4

   PIN FE_OFN10987_a_0_6_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 244.594 0.0 244.622 0.163 ;
      END
   END FE_OFN10987_a_0_6_1

   PIN FE_OFN10999_a_0_4_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 82.29 248.0 82.318 ;
      END
   END FE_OFN10999_a_0_4_7

   PIN FE_OFN11007_a_0_4_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 234.546 0.0 234.574 0.163 ;
      END
   END FE_OFN11007_a_0_4_0

   PIN FE_OFN12751_n_142961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.578 154.717 126.606 154.88 ;
      END
   END FE_OFN12751_n_142961

   PIN FE_OFN12753_n_142961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.77 154.717 110.798 154.88 ;
      END
   END FE_OFN12753_n_142961

   PIN FE_OFN14480_n_112183
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 133.746 154.717 133.774 154.88 ;
      END
   END FE_OFN14480_n_112183

   PIN FE_OFN14491_n_112182
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.81 154.717 133.838 154.88 ;
      END
   END FE_OFN14491_n_112182

   PIN FE_OFN14493_n_112182
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.578 154.717 150.606 154.88 ;
      END
   END FE_OFN14493_n_112182

   PIN FE_OFN14699_a_9_6_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 120.626 248.0 120.654 ;
      END
   END FE_OFN14699_a_9_6_7

   PIN FE_OFN14911_n_142849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.73 154.717 95.758 154.88 ;
      END
   END FE_OFN14911_n_142849

   PIN FE_OFN15367_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 140.658 248.0 140.686 ;
      END
   END FE_OFN15367_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_13_

   PIN FE_OFN15376_n_21671
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 53.042 248.0 53.07 ;
      END
   END FE_OFN15376_n_21671

   PIN FE_OFN15983_n_36821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.57 154.717 83.598 154.88 ;
      END
   END FE_OFN15983_n_36821

   PIN FE_OFN16026_a_0_6_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 242.546 0.0 242.574 0.163 ;
      END
   END FE_OFN16026_a_0_6_1

   PIN FE_OFN16151_a_2_4_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.322 0.0 238.35 0.163 ;
      END
   END FE_OFN16151_a_2_4_5

   PIN FE_OFN16443_a_7_4_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 82.354 248.0 82.382 ;
      END
   END FE_OFN16443_a_7_4_5

   PIN FE_OFN16476_a_2_6_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 7.154 248.0 7.182 ;
      END
   END FE_OFN16476_a_2_6_1

   PIN FE_OFN17481_n_126984
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.802 0.0 106.83 0.163 ;
      END
   END FE_OFN17481_n_126984

   PIN FE_OFN17555_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.162 154.717 122.19 154.88 ;
      END
   END FE_OFN17555_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_

   PIN FE_OFN18498_n_22234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 111.346 248.0 111.374 ;
      END
   END FE_OFN18498_n_22234

   PIN FE_OFN18638_a_7_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.762 0.0 235.79 0.163 ;
      END
   END FE_OFN18638_a_7_6_4

   PIN FE_OFN18656_a_3_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 243.058 0.0 243.086 0.163 ;
      END
   END FE_OFN18656_a_3_6_4

   PIN FE_OFN18679_a_1_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 229.81 0.0 229.838 0.163 ;
      END
   END FE_OFN18679_a_1_6_4

   PIN FE_OFN19318_a_8_8_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 140.722 248.0 140.75 ;
      END
   END FE_OFN19318_a_8_8_4

   PIN FE_OFN19321_a_4_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 222.322 0.0 222.35 0.163 ;
      END
   END FE_OFN19321_a_4_6_4

   PIN FE_OFN437_n_21145
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 49.202 248.0 49.23 ;
      END
   END FE_OFN437_n_21145

   PIN FE_OFN4661_n_142849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.082 154.717 76.11 154.88 ;
      END
   END FE_OFN4661_n_142849

   PIN FE_OFN4678_n_112357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.674 154.717 106.702 154.88 ;
      END
   END FE_OFN4678_n_112357

   PIN FE_OFN4703_n_143619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.058 154.717 99.086 154.88 ;
      END
   END FE_OFN4703_n_143619

   PIN FE_OFN4840_n_140222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.442 154.717 91.47 154.88 ;
      END
   END FE_OFN4840_n_140222

   PIN FE_OFN4981_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 247.837 150.386 248.0 150.414 ;
      END
   END FE_OFN4981_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_11_

   PIN FE_OFN4983_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 150.066 248.0 150.094 ;
      END
   END FE_OFN4983_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_10_

   PIN FE_OFN5000_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.122 154.717 195.15 154.88 ;
      END
   END FE_OFN5000_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_11_

   PIN FE_OFN636_n_11194
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.93 0.0 242.958 0.163 ;
      END
   END FE_OFN636_n_11194

   PIN FE_OFN638_n_8336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 4.85 248.0 4.878 ;
      END
   END FE_OFN638_n_8336

   PIN FE_OFN651_n_7003
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 22.13 248.0 22.158 ;
      END
   END FE_OFN651_n_7003

   PIN FE_OFN741_n_22817
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 156.786 0.0 156.814 0.163 ;
      END
   END FE_OFN741_n_22817

   PIN FE_OFN8951_n_6635
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 214.45 154.717 214.478 154.88 ;
      END
   END FE_OFN8951_n_6635

   PIN FE_OFN9215_delay_add_ln34_unr2_unr8_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 22.194 248.0 22.222 ;
      END
   END FE_OFN9215_delay_add_ln34_unr2_unr8_stage2_stallmux_q_13_

   PIN FE_OFN9217_delay_add_ln34_unr2_unr8_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 72.818 248.0 72.846 ;
      END
   END FE_OFN9217_delay_add_ln34_unr2_unr8_stage2_stallmux_q_12_

   PIN FE_OFN9884_b_4_8_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.082 154.717 4.11 154.88 ;
      END
   END FE_OFN9884_b_4_8_1

   PIN FE_OFN9902_b_4_7_9
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.082 154.717 84.11 154.88 ;
      END
   END FE_OFN9902_b_4_7_9

   PIN delay_add_ln34_unr2_unr1_stage2_stallmux_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 4.914 248.0 4.942 ;
      END
   END delay_add_ln34_unr2_unr1_stage2_stallmux_q_10_

   PIN delay_add_ln34_unr2_unr1_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 14.386 248.0 14.414 ;
      END
   END delay_add_ln34_unr2_unr1_stage2_stallmux_q_7_

   PIN delay_add_ln34_unr2_unr2_stage2_stallmux_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 101.618 248.0 101.646 ;
      END
   END delay_add_ln34_unr2_unr2_stage2_stallmux_q_1_

   PIN delay_add_ln34_unr2_unr2_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 7.09 248.0 7.118 ;
      END
   END delay_add_ln34_unr2_unr2_stage2_stallmux_q_2_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 206.77 0.0 206.798 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_12_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 202.866 0.0 202.894 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_14_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.21 0.0 172.238 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_7_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.69 0.0 160.718 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr3_unr7_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.898 154.717 102.926 154.88 ;
      END
   END delay_mul_ln34_unr3_unr7_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.514 154.717 166.542 154.88 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr4_unr7_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 187.442 0.0 187.47 0.163 ;
      END
   END delay_mul_ln34_unr4_unr7_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr4_unr9_stage2_stallmux_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 18.482 248.0 18.51 ;
      END
   END delay_mul_ln34_unr4_unr9_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 133.746 248.0 133.774 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.026 154.717 199.054 154.88 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.186 154.717 195.214 154.88 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 183.666 154.717 183.694 154.88 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 168.242 154.717 168.27 154.88 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.626 154.717 160.654 154.88 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_9_

   PIN mul_4646_72_n_150
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.706 154.717 110.734 154.88 ;
      END
   END mul_4646_72_n_150

   PIN mul_4646_72_n_251
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.994 154.717 107.022 154.88 ;
      END
   END mul_4646_72_n_251

   PIN mul_4646_72_n_58
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.546 0.0 114.574 0.163 ;
      END
   END mul_4646_72_n_58

   PIN mul_4646_72_n_59
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.426 0.0 125.454 0.163 ;
      END
   END mul_4646_72_n_59

   PIN mul_4646_72_n_75
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.594 0.0 124.622 0.163 ;
      END
   END mul_4646_72_n_75

   PIN mul_4646_72_n_756
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.45 0.0 134.478 0.163 ;
      END
   END mul_4646_72_n_756

   PIN mul_4650_72_n_212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.738 154.717 130.766 154.88 ;
      END
   END mul_4650_72_n_212

   PIN mul_4650_72_n_213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.354 154.717 130.382 154.88 ;
      END
   END mul_4650_72_n_213

   PIN mul_4650_72_n_214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.802 154.717 130.83 154.88 ;
      END
   END mul_4650_72_n_214

   PIN mul_4650_72_n_217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.362 0.0 45.39 0.163 ;
      END
   END mul_4650_72_n_217

   PIN mul_4650_72_n_239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.29 154.717 90.318 154.88 ;
      END
   END mul_4650_72_n_239

   PIN mul_4650_72_n_252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.554 154.717 37.582 154.88 ;
      END
   END mul_4650_72_n_252

   PIN mul_4650_72_n_285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.714 154.717 41.742 154.88 ;
      END
   END mul_4650_72_n_285

   PIN mul_4650_72_n_287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.65 154.717 41.678 154.88 ;
      END
   END mul_4650_72_n_287

   PIN mul_4650_72_n_289
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.858 154.717 55.886 154.88 ;
      END
   END mul_4650_72_n_289

   PIN mul_4650_72_n_292
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.002 154.717 30.03 154.88 ;
      END
   END mul_4650_72_n_292

   PIN mul_4650_72_n_311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.146 154.717 76.174 154.88 ;
      END
   END mul_4650_72_n_311

   PIN mul_4650_72_n_313
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.954 154.717 75.982 154.88 ;
      END
   END mul_4650_72_n_313

   PIN mul_4650_72_n_55
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.114 0.0 56.142 0.163 ;
      END
   END mul_4650_72_n_55

   PIN mul_4650_72_n_73
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.37 0.0 112.398 0.163 ;
      END
   END mul_4650_72_n_73

   PIN mul_4650_72_n_777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.234 0.0 53.262 0.163 ;
      END
   END mul_4650_72_n_777

   PIN mul_4650_72_n_78
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.682 154.717 133.71 154.88 ;
      END
   END mul_4650_72_n_78

   PIN mul_4650_72_n_848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.426 0.0 45.454 0.163 ;
      END
   END mul_4650_72_n_848

   PIN n_111907
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.082 154.717 148.11 154.88 ;
      END
   END n_111907

   PIN n_112284
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.906 154.717 33.934 154.88 ;
      END
   END n_112284

   PIN n_112720
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.258 154.717 126.286 154.88 ;
      END
   END n_112720

   PIN n_113639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.058 154.717 51.086 154.88 ;
      END
   END n_113639

   PIN n_113790
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.482 154.717 82.51 154.88 ;
      END
   END n_113790

   PIN n_114086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 118.45 154.717 118.478 154.88 ;
      END
   END n_114086

   PIN n_114387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.41 0.0 95.438 0.163 ;
      END
   END n_114387

   PIN n_114392
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.354 154.717 50.382 154.88 ;
      END
   END n_114392

   PIN n_114607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.77 0.0 94.798 0.163 ;
      END
   END n_114607

   PIN n_114644
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.242 154.717 120.27 154.88 ;
      END
   END n_114644

   PIN n_114654
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 68.53 154.717 68.558 154.88 ;
      END
   END n_114654

   PIN n_115067
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.146 0.0 76.174 0.163 ;
      END
   END n_115067

   PIN n_115075
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.946 154.717 56.974 154.88 ;
      END
   END n_115075

   PIN n_115173
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 57.01 154.717 57.038 154.88 ;
      END
   END n_115173

   PIN n_115193
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.642 154.717 110.67 154.88 ;
      END
   END n_115193

   PIN n_115538
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.642 154.717 118.67 154.88 ;
      END
   END n_115538

   PIN n_115592
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.466 154.717 68.494 154.88 ;
      END
   END n_115592

   PIN n_115601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.746 154.717 93.774 154.88 ;
      END
   END n_115601

   PIN n_115610
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.61 154.717 114.638 154.88 ;
      END
   END n_115610

   PIN n_115697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.106 154.717 109.134 154.88 ;
      END
   END n_115697

   PIN n_115863
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.706 154.717 30.734 154.88 ;
      END
   END n_115863

   PIN n_115878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.17 154.717 53.198 154.88 ;
      END
   END n_115878

   PIN n_115897
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.418 154.717 34.446 154.88 ;
      END
   END n_115897

   PIN n_116017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.218 154.717 111.246 154.88 ;
      END
   END n_116017

   PIN n_116364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.362 154.717 101.39 154.88 ;
      END
   END n_116364

   PIN n_116388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.346 154.717 63.374 154.88 ;
      END
   END n_116388

   PIN n_116530
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 126.13 154.717 126.158 154.88 ;
      END
   END n_116530

   PIN n_116580
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.85 154.717 92.878 154.88 ;
      END
   END n_116580

   PIN n_116853
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.994 154.717 107.022 154.88 ;
      END
   END n_116853

   PIN n_116869
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.786 154.717 60.814 154.88 ;
      END
   END n_116869

   PIN n_117308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.194 0.0 46.222 0.163 ;
      END
   END n_117308

   PIN n_117932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.77 154.717 46.798 154.88 ;
      END
   END n_117932

   PIN n_118446
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.066 154.717 118.094 154.88 ;
      END
   END n_118446

   PIN n_118851
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.226 154.717 50.254 154.88 ;
      END
   END n_118851

   PIN n_118961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.69 154.717 96.718 154.88 ;
      END
   END n_118961

   PIN n_119042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.73 154.717 103.758 154.88 ;
      END
   END n_119042

   PIN n_119323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.034 154.717 98.062 154.88 ;
      END
   END n_119323

   PIN n_119415
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.506 154.717 107.534 154.88 ;
      END
   END n_119415

   PIN n_119457
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.666 154.717 87.694 154.88 ;
      END
   END n_119457

   PIN n_120207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.45 154.717 118.478 154.88 ;
      END
   END n_120207

   PIN n_120352
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.21 0.0 76.238 0.163 ;
      END
   END n_120352

   PIN n_120375
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.546 154.717 114.574 154.88 ;
      END
   END n_120375

   PIN n_120599
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.994 0.0 107.022 0.163 ;
      END
   END n_120599

   PIN n_120600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.93 0.0 106.958 0.163 ;
      END
   END n_120600

   PIN n_121035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.002 154.717 118.03 154.88 ;
      END
   END n_121035

   PIN n_121273
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.13 0.0 46.158 0.163 ;
      END
   END n_121273

   PIN n_121548
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.266 154.717 17.294 154.88 ;
      END
   END n_121548

   PIN n_121555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.738 154.717 106.766 154.88 ;
      END
   END n_121555

   PIN n_121639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.674 154.717 114.702 154.88 ;
      END
   END n_121639

   PIN n_121887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.73 0.0 63.758 0.163 ;
      END
   END n_121887

   PIN n_121951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.722 0.0 92.75 0.163 ;
      END
   END n_121951

   PIN n_122050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.418 0.0 98.446 0.163 ;
      END
   END n_122050

   PIN n_122090
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.882 154.717 56.91 154.88 ;
      END
   END n_122090

   PIN n_122254
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.33 0.0 49.358 0.163 ;
      END
   END n_122254

   PIN n_122427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 110.962 0.163 110.99 ;
      END
   END n_122427

   PIN n_124381
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 95.346 0.163 95.374 ;
      END
   END n_124381

   PIN n_124384
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 87.666 0.163 87.694 ;
      END
   END n_124384

   PIN n_124473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.466 0.163 68.494 ;
      END
   END n_124473

   PIN n_124480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.226 154.717 26.254 154.88 ;
      END
   END n_124480

   PIN n_124768
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.61 154.717 138.638 154.88 ;
      END
   END n_124768

   PIN n_124884
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.946 154.717 128.974 154.88 ;
      END
   END n_124884

   PIN n_124890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.226 154.717 122.254 154.88 ;
      END
   END n_124890

   PIN n_124892
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.866 0.0 106.894 0.163 ;
      END
   END n_124892

   PIN n_125201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 91.762 0.163 91.79 ;
      END
   END n_125201

   PIN n_125438
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 133.81 0.0 133.838 0.163 ;
      END
   END n_125438

   PIN n_125484
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.65 0.0 89.678 0.163 ;
      END
   END n_125484

   PIN n_126152
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 91.442 0.163 91.47 ;
      END
   END n_126152

   PIN n_126230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 95.282 0.163 95.31 ;
      END
   END n_126230

   PIN n_126465
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.29 0.0 122.318 0.163 ;
      END
   END n_126465

   PIN n_126950
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.13 154.717 30.158 154.88 ;
      END
   END n_126950

   PIN n_127100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.074 0.0 65.102 0.163 ;
      END
   END n_127100

   PIN n_127101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.138 0.0 65.166 0.163 ;
      END
   END n_127101

   PIN n_127102
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.562 0.0 64.59 0.163 ;
      END
   END n_127102

   PIN n_127132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.418 154.717 122.446 154.88 ;
      END
   END n_127132

   PIN n_127133
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.354 154.717 122.382 154.88 ;
      END
   END n_127133

   PIN n_127136
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.93 0.0 106.958 0.163 ;
      END
   END n_127136

   PIN n_127563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.97 0.0 129.998 0.163 ;
      END
   END n_127563

   PIN n_128225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.09 0.0 7.118 0.163 ;
      END
   END n_128225

   PIN n_129278
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.586 0.0 41.614 0.163 ;
      END
   END n_129278

   PIN n_130041
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.714 0.0 41.742 0.163 ;
      END
   END n_130041

   PIN n_130821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 83.762 0.163 83.79 ;
      END
   END n_130821

   PIN n_131531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.546 0.163 114.574 ;
      END
   END n_131531

   PIN n_133774
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.682 0.0 61.71 0.163 ;
      END
   END n_133774

   PIN n_13498
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.882 154.717 152.91 154.88 ;
      END
   END n_13498

   PIN n_137441
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.378 0.0 139.406 0.163 ;
      END
   END n_137441

   PIN n_142793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.586 154.717 137.614 154.88 ;
      END
   END n_142793

   PIN n_142961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 95.346 248.0 95.374 ;
      END
   END n_142961

   PIN n_143003
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.826 154.717 83.854 154.88 ;
      END
   END n_143003

   PIN n_14932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.41 154.717 191.438 154.88 ;
      END
   END n_14932

   PIN n_14933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 188.85 154.717 188.878 154.88 ;
      END
   END n_14933

   PIN n_14966
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 190.194 154.717 190.222 154.88 ;
      END
   END n_14966

   PIN n_16625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 79.986 248.0 80.014 ;
      END
   END n_16625

   PIN n_16626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 80.114 248.0 80.142 ;
      END
   END n_16626

   PIN n_17619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 114.482 248.0 114.51 ;
      END
   END n_17619

   PIN n_19300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.794 154.717 159.822 154.88 ;
      END
   END n_19300

   PIN n_19852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.146 154.717 196.174 154.88 ;
      END
   END n_19852

   PIN n_19853
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.346 154.717 191.374 154.88 ;
      END
   END n_19853

   PIN n_20189
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 14.578 248.0 14.606 ;
      END
   END n_20189

   PIN n_20626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.338 154.717 164.366 154.88 ;
      END
   END n_20626

   PIN n_21390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 79.858 248.0 79.886 ;
      END
   END n_21390

   PIN n_21391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 82.418 248.0 82.446 ;
      END
   END n_21391

   PIN n_21448
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.69 154.717 160.718 154.88 ;
      END
   END n_21448

   PIN n_21461
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.314 0.0 203.342 0.163 ;
      END
   END n_21461

   PIN n_21505
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 150.13 248.0 150.158 ;
      END
   END n_21505

   PIN n_21517
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 137.522 248.0 137.55 ;
      END
   END n_21517

   PIN n_21590
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 168.37 154.717 168.398 154.88 ;
      END
   END n_21590

   PIN n_21591
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 168.306 154.717 168.334 154.88 ;
      END
   END n_21591

   PIN n_21678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 183.73 154.717 183.758 154.88 ;
      END
   END n_21678

   PIN n_21692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 247.837 150.45 248.0 150.478 ;
      END
   END n_21692

   PIN n_21696
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 72.882 248.0 72.91 ;
      END
   END n_21696

   PIN n_21711
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 137.586 248.0 137.614 ;
      END
   END n_21711

   PIN n_21955
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.106 0.0 149.134 0.163 ;
      END
   END n_21955

   PIN n_21973
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 80.05 248.0 80.078 ;
      END
   END n_21973

   PIN n_21974
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 79.922 248.0 79.95 ;
      END
   END n_21974

   PIN n_21990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 29.938 248.0 29.966 ;
      END
   END n_21990

   PIN n_22100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.042 0.0 149.07 0.163 ;
      END
   END n_22100

   PIN n_22130
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 150.322 248.0 150.35 ;
      END
   END n_22130

   PIN n_22131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 145.202 248.0 145.23 ;
      END
   END n_22131

   PIN n_22132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 150.194 248.0 150.222 ;
      END
   END n_22132

   PIN n_22135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 72.562 248.0 72.59 ;
      END
   END n_22135

   PIN n_22222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 187.57 154.717 187.598 154.88 ;
      END
   END n_22222

   PIN n_22223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 160.69 154.717 160.718 154.88 ;
      END
   END n_22223

   PIN n_22241
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 114.546 248.0 114.574 ;
      END
   END n_22241

   PIN n_22502
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 168.37 0.0 168.398 0.163 ;
      END
   END n_22502

   PIN n_22542
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 34.418 248.0 34.446 ;
      END
   END n_22542

   PIN n_23096
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 23.922 248.0 23.95 ;
      END
   END n_23096

   PIN n_23324
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 68.466 248.0 68.494 ;
      END
   END n_23324

   PIN n_23325
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 91.25 248.0 91.278 ;
      END
   END n_23325

   PIN n_23968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 122.098 248.0 122.126 ;
      END
   END n_23968

   PIN n_23969
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 118.386 248.0 118.414 ;
      END
   END n_23969

   PIN n_23973
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 120.69 248.0 120.718 ;
      END
   END n_23973

   PIN n_24209
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.042 154.717 149.07 154.88 ;
      END
   END n_24209

   PIN n_24210
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.01 154.717 129.038 154.88 ;
      END
   END n_24210

   PIN n_24293
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 87.602 248.0 87.63 ;
      END
   END n_24293

   PIN n_24393
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 76.146 248.0 76.174 ;
      END
   END n_24393

   PIN n_24834
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.994 154.717 155.022 154.88 ;
      END
   END n_24834

   PIN n_24836
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.482 154.717 154.51 154.88 ;
      END
   END n_24836

   PIN n_24845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.97 154.717 145.998 154.88 ;
      END
   END n_24845

   PIN n_24847
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.906 154.717 145.934 154.88 ;
      END
   END n_24847

   PIN n_24890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 133.81 248.0 133.838 ;
      END
   END n_24890

   PIN n_24892
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 137.65 248.0 137.678 ;
      END
   END n_24892

   PIN n_24997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 131.058 248.0 131.086 ;
      END
   END n_24997

   PIN n_25050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 210.61 154.717 210.638 154.88 ;
      END
   END n_25050

   PIN n_25074
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 153.01 154.717 153.038 154.88 ;
      END
   END n_25074

   PIN n_25101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 133.682 248.0 133.71 ;
      END
   END n_25101

   PIN n_25132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 92.018 248.0 92.046 ;
      END
   END n_25132

   PIN n_25257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.842 154.717 145.87 154.88 ;
      END
   END n_25257

   PIN n_25529
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 150.514 154.717 150.542 154.88 ;
      END
   END n_25529

   PIN n_25531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.106 154.717 149.134 154.88 ;
      END
   END n_25531

   PIN n_25624
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 92.082 248.0 92.11 ;
      END
   END n_25624

   PIN n_26550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 101.746 248.0 101.774 ;
      END
   END n_26550

   PIN n_26818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 101.682 248.0 101.71 ;
      END
   END n_26818

   PIN n_27649
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 233.65 154.717 233.678 154.88 ;
      END
   END n_27649

   PIN n_27650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.074 154.717 241.102 154.88 ;
      END
   END n_27650

   PIN n_27752
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.25 154.717 195.278 154.88 ;
      END
   END n_27752

   PIN n_2800
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.786 0.163 60.814 ;
      END
   END n_2800

   PIN n_28028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.746 154.717 229.774 154.88 ;
      END
   END n_28028

   PIN n_28030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.466 154.717 228.494 154.88 ;
      END
   END n_28030

   PIN n_28637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.786 154.717 180.814 154.88 ;
      END
   END n_28637

   PIN n_28704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 192.498 0.0 192.526 0.163 ;
      END
   END n_28704

   PIN n_28825
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 150.258 248.0 150.286 ;
      END
   END n_28825

   PIN n_29574
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 145.138 248.0 145.166 ;
      END
   END n_29574

   PIN n_29646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 140.786 248.0 140.814 ;
      END
   END n_29646

   PIN n_32056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.194 154.717 78.222 154.88 ;
      END
   END n_32056

   PIN n_32073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.986 154.717 88.014 154.88 ;
      END
   END n_32073

   PIN n_32468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.114 154.717 112.142 154.88 ;
      END
   END n_32468

   PIN n_32697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.426 0.163 101.454 ;
      END
   END n_32697

   PIN n_32704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.49 154.717 45.518 154.88 ;
      END
   END n_32704

   PIN n_32867
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.362 0.163 101.39 ;
      END
   END n_32867

   PIN n_33365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.49 0.163 101.518 ;
      END
   END n_33365

   PIN n_33776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 131.25 154.717 131.278 154.88 ;
      END
   END n_33776

   PIN n_34364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.402 154.717 60.43 154.88 ;
      END
   END n_34364

   PIN n_34374
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.978 154.717 53.006 154.88 ;
      END
   END n_34374

   PIN n_34614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.93 154.717 106.958 154.88 ;
      END
   END n_34614

   PIN n_34686
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 133.682 154.717 133.71 154.88 ;
      END
   END n_34686

   PIN n_35435
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.13 154.717 38.158 154.88 ;
      END
   END n_35435

   PIN n_35467
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.866 154.717 106.894 154.88 ;
      END
   END n_35467

   PIN n_36948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.53 154.717 68.558 154.88 ;
      END
   END n_36948

   PIN n_37020
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.49 154.717 69.518 154.88 ;
      END
   END n_37020

   PIN n_37253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.082 154.717 76.11 154.88 ;
      END
   END n_37253

   PIN n_37497
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.458 154.717 25.486 154.88 ;
      END
   END n_37497

   PIN n_37498
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.826 154.717 19.854 154.88 ;
      END
   END n_37498

   PIN n_37637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.474 154.717 95.502 154.88 ;
      END
   END n_37637

   PIN n_38077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.01 0.0 113.038 0.163 ;
      END
   END n_38077

   PIN n_39307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.026 0.0 103.054 0.163 ;
      END
   END n_39307

   PIN n_39821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 131.122 248.0 131.15 ;
      END
   END n_39821

   PIN n_39967
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 44.018 248.0 44.046 ;
      END
   END n_39967

   PIN n_40268
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 23.986 248.0 24.014 ;
      END
   END n_40268

   PIN n_40473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.69 0.0 208.718 0.163 ;
      END
   END n_40473

   PIN n_40638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.602 0.0 239.63 0.163 ;
      END
   END n_40638

   PIN n_40714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 83.634 248.0 83.662 ;
      END
   END n_40714

   PIN n_41448
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.266 154.717 145.294 154.88 ;
      END
   END n_41448

   PIN n_44877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.026 154.717 103.054 154.88 ;
      END
   END n_44877

   PIN n_47745
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.698 154.717 83.726 154.88 ;
      END
   END n_47745

   PIN n_47887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.146 154.717 76.174 154.88 ;
      END
   END n_47887

   PIN n_48179
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.97 154.717 73.998 154.88 ;
      END
   END n_48179

   PIN n_54122
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.65 154.717 41.678 154.88 ;
      END
   END n_54122

   PIN n_54294
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.402 154.717 68.43 154.88 ;
      END
   END n_54294

   PIN n_5456
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.866 0.0 106.894 0.163 ;
      END
   END n_5456

   PIN n_5457
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.706 0.0 110.734 0.163 ;
      END
   END n_5457

   PIN n_57601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.434 154.717 72.462 154.88 ;
      END
   END n_57601

   PIN n_59902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.834 154.717 54.862 154.88 ;
      END
   END n_59902

   PIN n_60533
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.306 154.717 72.334 154.88 ;
      END
   END n_60533

   PIN n_62170
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.018 154.717 76.046 154.88 ;
      END
   END n_62170

   PIN n_6519
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 237.49 154.717 237.518 154.88 ;
      END
   END n_6519

   PIN n_65559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 219.442 0.0 219.47 0.163 ;
      END
   END n_65559

   PIN n_7333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 6.962 248.0 6.99 ;
      END
   END n_7333

   PIN n_8253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.386 0.0 150.414 0.163 ;
      END
   END n_8253

   PIN n_9777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 247.837 79.986 248.0 80.014 ;
      END
   END n_9777

   PIN FE_OCPN15632_n_40178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.378 0.0 211.406 0.163 ;
      END
   END FE_OCPN15632_n_40178

   PIN FE_OFN10061_b_4_3_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.354 154.717 74.382 154.88 ;
      END
   END FE_OFN10061_b_4_3_6

   PIN FE_OFN10064_b_4_3_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.578 154.717 110.606 154.88 ;
      END
   END FE_OFN10064_b_4_3_5

   PIN FE_OFN10067_b_4_3_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.338 154.717 92.366 154.88 ;
      END
   END FE_OFN10067_b_4_3_4

   PIN FE_OFN10070_b_4_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.41 154.717 95.438 154.88 ;
      END
   END FE_OFN10070_b_4_3_3

   PIN FE_OFN10072_b_4_3_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.546 154.717 114.574 154.88 ;
      END
   END FE_OFN10072_b_4_3_2

   PIN FE_OFN10076_b_4_3_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.506 154.717 91.534 154.88 ;
      END
   END FE_OFN10076_b_4_3_1

   PIN FE_OFN10077_b_4_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.378 154.717 91.406 154.88 ;
      END
   END FE_OFN10077_b_4_3_0

   PIN FE_OFN10078_b_4_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.25 154.717 99.278 154.88 ;
      END
   END FE_OFN10078_b_4_3_0

   PIN FE_OFN10180_b_4_0_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.65 154.798 65.678 154.88 ;
      END
   END FE_OFN10180_b_4_0_3

   PIN FE_OFN10188_b_4_0_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.066 154.717 126.094 154.88 ;
      END
   END FE_OFN10188_b_4_0_0

   PIN FE_OFN10818_a_3_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 202.93 154.717 202.958 154.88 ;
      END
   END FE_OFN10818_a_3_6_7

   PIN FE_OFN10857_a_2_8_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 244.978 154.717 245.006 154.88 ;
      END
   END FE_OFN10857_a_2_8_1

   PIN FE_OFN10871_a_2_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.29 154.717 218.318 154.88 ;
      END
   END FE_OFN10871_a_2_6_7

   PIN FE_OFN10986_a_0_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 240.69 154.717 240.718 154.88 ;
      END
   END FE_OFN10986_a_0_6_1

   PIN FE_OFN11519_n_40714
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 83.698 248.0 83.726 ;
      END
   END FE_OFN11519_n_40714

   PIN FE_OFN11549_n_142793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.842 154.717 113.87 154.88 ;
      END
   END FE_OFN11549_n_142793

   PIN FE_OFN1154_n_10378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.33 0.0 145.358 0.163 ;
      END
   END FE_OFN1154_n_10378

   PIN FE_OFN11610_n_39244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.002 154.717 126.03 154.88 ;
      END
   END FE_OFN11610_n_39244

   PIN FE_OFN11880_n_143202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.378 154.717 99.406 154.88 ;
      END
   END FE_OFN11880_n_143202

   PIN FE_OFN11883_n_143200
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.474 154.717 87.502 154.88 ;
      END
   END FE_OFN11883_n_143200

   PIN FE_OFN12031_n_143507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.826 154.717 83.854 154.88 ;
      END
   END FE_OFN12031_n_143507

   PIN FE_OFN12057_n_140222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 187.506 154.717 187.534 154.88 ;
      END
   END FE_OFN12057_n_140222

   PIN FE_OFN12086_n_143619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.946 154.717 96.974 154.88 ;
      END
   END FE_OFN12086_n_143619

   PIN FE_OFN12427_n_143003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.482 154.717 82.51 154.88 ;
      END
   END FE_OFN12427_n_143003

   PIN FE_OFN12759_n_142961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.314 154.717 99.342 154.88 ;
      END
   END FE_OFN12759_n_142961

   PIN FE_OFN13003_n_39130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.314 154.717 99.342 154.88 ;
      END
   END FE_OFN13003_n_39130

   PIN FE_OFN13192_n_37615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.41 154.717 87.438 154.88 ;
      END
   END FE_OFN13192_n_37615

   PIN FE_OFN13223_n_143620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.826 154.717 99.854 154.88 ;
      END
   END FE_OFN13223_n_143620

   PIN FE_OFN13288_n_143034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.242 154.717 96.27 154.88 ;
      END
   END FE_OFN13288_n_143034

   PIN FE_OFN13294_n_143033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.018 154.717 84.046 154.88 ;
      END
   END FE_OFN13294_n_143033

   PIN FE_OFN13296_n_143032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.954 154.717 91.982 154.88 ;
      END
   END FE_OFN13296_n_143032

   PIN FE_OFN13353_n_142795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.778 154.717 113.806 154.88 ;
      END
   END FE_OFN13353_n_142795

   PIN FE_OFN13512_n_112357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.618 154.717 77.646 154.88 ;
      END
   END FE_OFN13512_n_112357

   PIN FE_OFN13586_n_143006
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.97 154.717 89.998 154.88 ;
      END
   END FE_OFN13586_n_143006

   PIN FE_OFN14074_n_142964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.154 154.717 95.182 154.88 ;
      END
   END FE_OFN14074_n_142964

   PIN FE_OFN14079_n_142963
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.05 154.717 88.078 154.88 ;
      END
   END FE_OFN14079_n_142963

   PIN FE_OFN14083_n_142962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.338 154.717 68.366 154.88 ;
      END
   END FE_OFN14083_n_142962

   PIN FE_OFN14327_n_140207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.186 154.798 91.214 154.88 ;
      END
   END FE_OFN14327_n_140207

   PIN FE_OFN14360_n_143300
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.106 154.717 53.134 154.88 ;
      END
   END FE_OFN14360_n_143300

   PIN FE_OFN14403_n_142794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.05 154.717 88.078 154.88 ;
      END
   END FE_OFN14403_n_142794

   PIN FE_OFN14479_n_112183
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.794 154.717 143.822 154.88 ;
      END
   END FE_OFN14479_n_112183

   PIN FE_OFN14487_n_143005
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.706 154.717 102.734 154.88 ;
      END
   END FE_OFN14487_n_143005

   PIN FE_OFN14698_a_9_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 202.866 154.717 202.894 154.88 ;
      END
   END FE_OFN14698_a_9_6_7

   PIN FE_OFN14912_n_142849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.282 154.717 95.31 154.88 ;
      END
   END FE_OFN14912_n_142849

   PIN FE_OFN14984_n_112030
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.434 154.717 128.462 154.88 ;
      END
   END FE_OFN14984_n_112030

   PIN FE_OFN15130_n_20599
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 247.026 0.0 247.054 0.163 ;
      END
   END FE_OFN15130_n_20599

   PIN FE_OFN15291_n_111917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.186 154.717 99.214 154.88 ;
      END
   END FE_OFN15291_n_111917

   PIN FE_OFN15295_n_111917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.482 154.717 114.51 154.88 ;
      END
   END FE_OFN15295_n_111917

   PIN FE_OFN15366_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.018 0.0 212.046 0.163 ;
      END
   END FE_OFN15366_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_13_

   PIN FE_OFN15383_n_22225
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 240.434 0.0 240.462 0.163 ;
      END
   END FE_OFN15383_n_22225

   PIN FE_OFN15982_n_36821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.538 154.717 79.566 154.88 ;
      END
   END FE_OFN15982_n_36821

   PIN FE_OFN16234_n_40172
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 43.954 248.0 43.982 ;
      END
   END FE_OFN16234_n_40172

   PIN FE_OFN16237_n_40170
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.69 0.0 224.718 0.163 ;
      END
   END FE_OFN16237_n_40170

   PIN FE_OFN16239_n_40166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.682 0.0 229.71 0.163 ;
      END
   END FE_OFN16239_n_40166

   PIN FE_OFN16241_n_40166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 43.89 248.0 43.918 ;
      END
   END FE_OFN16241_n_40166

   PIN FE_OFN16256_n_40159
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 235.25 0.0 235.278 0.163 ;
      END
   END FE_OFN16256_n_40159

   PIN FE_OFN16649_n_7003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 26.226 248.0 26.254 ;
      END
   END FE_OFN16649_n_7003

   PIN FE_OFN17473_n_142961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 106.866 248.0 106.894 ;
      END
   END FE_OFN17473_n_142961

   PIN FE_OFN17490_n_142849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.802 154.717 106.83 154.88 ;
      END
   END FE_OFN17490_n_142849

   PIN FE_OFN17556_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.29 154.717 122.318 154.88 ;
      END
   END FE_OFN17556_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_

   PIN FE_OFN18570_b_4_7_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.706 154.717 14.734 154.88 ;
      END
   END FE_OFN18570_b_4_7_9

   PIN FE_OFN4555_n_142963
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.178 154.717 72.206 154.88 ;
      END
   END FE_OFN4555_n_142963

   PIN FE_OFN4568_n_41387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.978 154.717 149.006 154.88 ;
      END
   END FE_OFN4568_n_41387

   PIN FE_OFN4613_n_142796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 87.602 154.717 87.63 154.88 ;
      END
   END FE_OFN4613_n_142796

   PIN FE_OFN4646_n_142850
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.778 154.798 65.806 154.88 ;
      END
   END FE_OFN4646_n_142850

   PIN FE_OFN4665_n_137232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.898 154.717 86.926 154.88 ;
      END
   END FE_OFN4665_n_137232

   PIN FE_OFN4702_n_143619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 87.73 154.717 87.758 154.88 ;
      END
   END FE_OFN4702_n_143619

   PIN FE_OFN4762_n_137230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.178 154.717 80.206 154.88 ;
      END
   END FE_OFN4762_n_137230

   PIN FE_OFN4773_n_143004
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.09 154.717 103.118 154.88 ;
      END
   END FE_OFN4773_n_143004

   PIN FE_OFN4784_n_143003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.61 154.717 18.638 154.88 ;
      END
   END FE_OFN4784_n_143003

   PIN FE_OFN4791_n_41686
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.026 154.717 103.054 154.88 ;
      END
   END FE_OFN4791_n_41686

   PIN FE_OFN4796_n_143145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.938 154.717 93.966 154.88 ;
      END
   END FE_OFN4796_n_143145

   PIN FE_OFN4798_n_143146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.938 154.717 93.966 154.88 ;
      END
   END FE_OFN4798_n_143146

   PIN FE_OFN4806_n_143143
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.122 154.717 99.15 154.88 ;
      END
   END FE_OFN4806_n_143143

   PIN FE_OFN4826_n_143199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.562 154.717 64.59 154.88 ;
      END
   END FE_OFN4826_n_143199

   PIN FE_OFN4885_n_36821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.986 154.717 80.014 154.88 ;
      END
   END FE_OFN4885_n_36821

   PIN FE_OFN4999_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 22.258 248.0 22.286 ;
      END
   END FE_OFN4999_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_11_

   PIN FE_OFN635_n_11194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.994 0.0 243.022 0.163 ;
      END
   END FE_OFN635_n_11194

   PIN FE_OFN637_n_8336
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.234 0.0 245.262 0.163 ;
      END
   END FE_OFN637_n_8336

   PIN FE_OFN654_n_8338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 244.018 0.0 244.046 0.163 ;
      END
   END FE_OFN654_n_8338

   PIN FE_OFN747_n_22238
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.89 0.0 83.918 0.163 ;
      END
   END FE_OFN747_n_22238

   PIN FE_OFN7582_n_40036
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 229.746 0.0 229.774 0.163 ;
      END
   END FE_OFN7582_n_40036

   PIN FE_OFN758_n_21703
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.282 0.0 199.31 0.163 ;
      END
   END FE_OFN758_n_21703

   PIN FE_OFN7819_n_40176
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 218.546 0.0 218.574 0.163 ;
      END
   END FE_OFN7819_n_40176

   PIN FE_OFN9214_delay_add_ln34_unr2_unr8_stage2_stallmux_q_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 10.802 248.0 10.83 ;
      END
   END FE_OFN9214_delay_add_ln34_unr2_unr8_stage2_stallmux_q_13_

   PIN FE_OFN9216_delay_add_ln34_unr2_unr8_stage2_stallmux_q_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 72.754 248.0 72.782 ;
      END
   END FE_OFN9216_delay_add_ln34_unr2_unr8_stage2_stallmux_q_12_

   PIN FE_OFN9895_b_4_7_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.922 154.717 79.95 154.88 ;
      END
   END FE_OFN9895_b_4_7_12

   PIN FE_OFN9897_b_4_7_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 73.714 154.717 73.742 154.88 ;
      END
   END FE_OFN9897_b_4_7_11

   PIN FE_OFN9899_b_4_7_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.89 154.717 83.918 154.88 ;
      END
   END FE_OFN9899_b_4_7_10

   PIN FE_OFN9905_b_4_7_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.514 154.717 70.542 154.88 ;
      END
   END FE_OFN9905_b_4_7_8

   PIN FE_OFN9908_b_4_7_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.21 154.717 76.238 154.88 ;
      END
   END FE_OFN9908_b_4_7_7

   PIN FE_OFN9910_b_4_7_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 80.05 154.717 80.078 154.88 ;
      END
   END FE_OFN9910_b_4_7_6

   PIN FE_OFN9911_b_4_7_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.242 154.717 72.27 154.88 ;
      END
   END FE_OFN9911_b_4_7_6

   PIN FE_OFN9913_b_4_7_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.858 154.717 87.886 154.88 ;
      END
   END FE_OFN9913_b_4_7_5

   PIN FE_OFN9914_b_4_7_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.866 154.717 106.894 154.88 ;
      END
   END FE_OFN9914_b_4_7_5

   PIN FE_OFN9916_b_4_7_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.89 154.717 83.918 154.88 ;
      END
   END FE_OFN9916_b_4_7_4

   PIN FE_OFN9917_b_4_7_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.57 154.717 99.598 154.88 ;
      END
   END FE_OFN9917_b_4_7_4

   PIN FE_OFN9919_b_4_7_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.954 154.717 83.982 154.88 ;
      END
   END FE_OFN9919_b_4_7_3

   PIN FE_OFN9920_b_4_7_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.442 154.717 91.47 154.88 ;
      END
   END FE_OFN9920_b_4_7_3

   PIN FE_OFN9922_b_4_7_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.538 154.717 87.566 154.88 ;
      END
   END FE_OFN9922_b_4_7_2

   PIN FE_OFN9923_b_4_7_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.482 154.717 106.51 154.88 ;
      END
   END FE_OFN9923_b_4_7_2

   PIN FE_OFN9925_b_4_7_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.93 154.717 50.958 154.88 ;
      END
   END FE_OFN9925_b_4_7_1

   PIN FE_OFN9928_b_4_7_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.722 154.717 76.75 154.88 ;
      END
   END FE_OFN9928_b_4_7_0

   PIN a_0_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 82.226 248.0 82.254 ;
      END
   END a_0_4_0

   PIN a_0_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 101.426 248.0 101.454 ;
      END
   END a_0_4_7

   PIN a_0_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 145.266 0.163 145.294 ;
      END
   END a_0_6_4

   PIN a_1_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 106.866 0.163 106.894 ;
      END
   END a_1_4_0

   PIN a_1_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 237.682 0.0 237.71 0.163 ;
      END
   END a_1_4_1

   PIN a_1_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 215.282 0.0 215.31 0.163 ;
      END
   END a_1_4_6

   PIN a_1_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.562 0.163 72.59 ;
      END
   END a_1_6_1

   PIN a_1_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 219.058 154.717 219.086 154.88 ;
      END
   END a_1_6_4

   PIN a_2_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 111.09 248.0 111.118 ;
      END
   END a_2_4_0

   PIN a_2_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.762 0.163 43.79 ;
      END
   END a_2_4_1

   PIN a_2_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 99.186 0.163 99.214 ;
      END
   END a_2_4_5

   PIN a_2_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 111.026 248.0 111.054 ;
      END
   END a_2_4_7

   PIN a_2_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 152.946 0.163 152.974 ;
      END
   END a_2_6_1

   PIN a_2_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 130.802 0.163 130.83 ;
      END
   END a_2_6_4

   PIN a_2_8_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 130.93 248.0 130.958 ;
      END
   END a_2_8_4

   PIN a_3_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 110.962 248.0 110.99 ;
      END
   END a_3_4_0

   PIN a_3_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.162 0.163 82.19 ;
      END
   END a_3_4_5

   PIN a_3_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.09 154.717 7.118 154.88 ;
      END
   END a_3_4_6

   PIN a_3_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.314 0.0 235.342 0.163 ;
      END
   END a_3_6_1

   PIN a_3_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 120.562 248.0 120.59 ;
      END
   END a_3_6_4

   PIN a_3_8_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 130.866 248.0 130.894 ;
      END
   END a_3_8_7

   PIN a_4_0_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 91.89 248.0 91.918 ;
      END
   END a_4_0_5

   PIN a_4_2_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 246.45 0.0 246.478 0.163 ;
      END
   END a_4_2_1

   PIN a_4_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.13 154.717 30.158 154.88 ;
      END
   END a_4_4_4

   PIN a_4_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 111.026 0.163 111.054 ;
      END
   END a_4_6_4

   PIN a_5_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.818 0.0 224.846 0.163 ;
      END
   END a_5_6_1

   PIN a_5_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 140.402 0.163 140.43 ;
      END
   END a_5_6_4

   PIN a_6_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.93 154.717 10.958 154.88 ;
      END
   END a_6_4_1

   PIN a_6_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.362 0.163 53.39 ;
      END
   END a_6_6_1

   PIN a_7_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.25 154.717 3.278 154.88 ;
      END
   END a_7_4_1

   PIN a_7_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 91.826 248.0 91.854 ;
      END
   END a_7_4_5

   PIN a_7_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.386 0.163 118.414 ;
      END
   END a_7_6_4

   PIN a_8_8_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 140.53 248.0 140.558 ;
      END
   END a_8_8_4

   PIN a_9_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 130.802 248.0 130.83 ;
      END
   END a_9_4_0

   PIN b_4_8_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 150.002 0.163 150.03 ;
      END
   END b_4_8_1

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.122 0.0 211.15 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_0_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 30.066 248.0 30.094 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_5_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 199.09 0.0 199.118 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_6_

   PIN delay_add_ln34_unr2_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 18.546 248.0 18.574 ;
      END
   END delay_add_ln34_unr2_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr3_unr0_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.298 0.0 157.326 0.163 ;
      END
   END delay_mul_ln34_unr3_unr0_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr3_unr5_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 242.482 0.0 242.51 0.163 ;
      END
   END delay_mul_ln34_unr3_unr5_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr3_unr7_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.866 0.0 218.894 0.163 ;
      END
   END delay_mul_ln34_unr3_unr7_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr3_unr7_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 34.29 248.0 34.318 ;
      END
   END delay_mul_ln34_unr3_unr7_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr3_unr7_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 194.93 0.0 194.958 0.163 ;
      END
   END delay_mul_ln34_unr3_unr7_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr3_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 53.426 248.0 53.454 ;
      END
   END delay_mul_ln34_unr3_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 63.154 248.0 63.182 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.65 154.717 137.678 154.88 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 141.49 154.717 141.518 154.88 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 184.498 154.717 184.526 154.88 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_z_7_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.762 154.717 83.79 154.88 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.946 154.717 56.974 154.88 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 206.706 0.0 206.734 0.163 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.466 0.0 220.494 0.163 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 210.546 0.0 210.574 0.163 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 140.466 248.0 140.494 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 217.01 0.0 217.038 0.163 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 10.93 248.0 10.958 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 37.81 248.0 37.838 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 41.522 248.0 41.55 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 37.746 248.0 37.774 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 41.586 248.0 41.614 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 87.73 248.0 87.758 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr5_unr5_stage2_stallmux_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 227.314 0.0 227.342 0.163 ;
      END
   END delay_mul_ln34_unr5_unr5_stage2_stallmux_z_10_

   PIN delay_mul_ln34_unr5_unr5_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.098 0.0 186.126 0.163 ;
      END
   END delay_mul_ln34_unr5_unr5_stage2_stallmux_z_11_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 140.402 248.0 140.43 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 26.29 248.0 26.318 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 126.13 0.0 126.158 0.163 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 181.042 0.0 181.07 0.163 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 60.786 248.0 60.814 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 3.186 248.0 3.214 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 7.026 248.0 7.054 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_8_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 3.122 248.0 3.15 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_9_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 133.874 154.798 133.902 154.88 ;
      END
   END ispd_clk

   PIN mul_4646_72_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.794 154.717 79.822 154.88 ;
      END
   END mul_4646_72_n_116

   PIN mul_4646_72_n_124
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.73 154.717 79.758 154.88 ;
      END
   END mul_4646_72_n_124

   PIN mul_4646_72_n_212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.218 154.717 95.246 154.88 ;
      END
   END mul_4646_72_n_212

   PIN mul_4646_72_n_213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.546 154.717 146.574 154.88 ;
      END
   END mul_4646_72_n_213

   PIN mul_4646_72_n_214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.13 154.717 126.158 154.88 ;
      END
   END mul_4646_72_n_214

   PIN mul_4646_72_n_96
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.794 154.717 87.822 154.88 ;
      END
   END mul_4646_72_n_96

   PIN mul_4646_72_n_97
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.426 0.0 101.454 0.163 ;
      END
   END mul_4646_72_n_97

   PIN mul_4646_72_n_98
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.49 0.0 101.518 0.163 ;
      END
   END mul_4646_72_n_98

   PIN mul_4650_72_n_288
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.482 154.717 58.51 154.88 ;
      END
   END mul_4650_72_n_288

   PIN mul_4650_72_n_307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.13 154.717 62.158 154.88 ;
      END
   END mul_4650_72_n_307

   PIN mul_4650_72_n_312
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.634 154.717 83.662 154.88 ;
      END
   END mul_4650_72_n_312

   PIN mul_4650_72_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.322 0.163 118.35 ;
      END
   END mul_4650_72_n_50

   PIN mul_4650_72_n_51
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.026 0.163 63.054 ;
      END
   END mul_4650_72_n_51

   PIN mul_4650_72_n_57
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.674 0.0 106.702 0.163 ;
      END
   END mul_4650_72_n_57

   PIN mul_4650_72_n_66
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.866 154.717 42.894 154.88 ;
      END
   END mul_4650_72_n_66

   PIN mul_4650_72_n_67
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.962 0.163 62.99 ;
      END
   END mul_4650_72_n_67

   PIN mul_4650_72_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.17 0.0 53.198 0.163 ;
      END
   END mul_4650_72_n_71

   PIN mul_4650_72_n_752
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.01 154.717 153.038 154.88 ;
      END
   END mul_4650_72_n_752

   PIN mul_4650_72_n_767
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.77 0.0 110.798 0.163 ;
      END
   END mul_4650_72_n_767

   PIN mul_4650_72_n_773
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.106 0.0 53.134 0.163 ;
      END
   END mul_4650_72_n_773

   PIN mul_4650_72_n_789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.562 0.163 64.59 ;
      END
   END mul_4650_72_n_789

   PIN mul_4650_72_n_837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.362 0.0 61.39 0.163 ;
      END
   END mul_4650_72_n_837

   PIN mul_4650_72_n_840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.65 0.0 41.678 0.163 ;
      END
   END mul_4650_72_n_840

   PIN n_112253
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.202 154.717 33.23 154.88 ;
      END
   END n_112253

   PIN n_112259
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.354 154.717 146.382 154.88 ;
      END
   END n_112259

   PIN n_112755
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.53 154.717 132.558 154.88 ;
      END
   END n_112755

   PIN n_113329
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.154 154.717 103.182 154.88 ;
      END
   END n_113329

   PIN n_113795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.09 154.717 103.118 154.88 ;
      END
   END n_113795

   PIN n_113875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.378 0.0 91.406 0.163 ;
      END
   END n_113875

   PIN n_114487
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.354 154.717 82.382 154.88 ;
      END
   END n_114487

   PIN n_115523
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.826 154.717 51.854 154.88 ;
      END
   END n_115523

   PIN n_115564
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.482 154.717 114.51 154.88 ;
      END
   END n_115564

   PIN n_115565
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.554 154.717 117.582 154.88 ;
      END
   END n_115565

   PIN n_116610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.898 154.717 46.926 154.88 ;
      END
   END n_116610

   PIN n_116849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.938 154.717 117.966 154.88 ;
      END
   END n_116849

   PIN n_116850
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.49 154.717 117.518 154.88 ;
      END
   END n_116850

   PIN n_117661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.962 154.717 102.99 154.88 ;
      END
   END n_117661

   PIN n_117721
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.346 0.0 95.374 0.163 ;
      END
   END n_117721

   PIN n_119045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.466 154.717 20.494 154.88 ;
      END
   END n_119045

   PIN n_120348
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.362 154.717 45.39 154.88 ;
      END
   END n_120348

   PIN n_120860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.042 154.717 53.07 154.88 ;
      END
   END n_120860

   PIN n_121613
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.178 154.717 24.206 154.88 ;
      END
   END n_121613

   PIN n_121641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 122.226 154.717 122.254 154.88 ;
      END
   END n_121641

   PIN n_121888
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.498 0.0 64.526 0.163 ;
      END
   END n_121888

   PIN n_123339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.426 154.717 45.454 154.88 ;
      END
   END n_123339

   PIN n_124376
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.794 0.0 63.822 0.163 ;
      END
   END n_124376

   PIN n_124377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.426 0.0 69.454 0.163 ;
      END
   END n_124377

   PIN n_124389
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.722 154.717 60.75 154.88 ;
      END
   END n_124389

   PIN n_124393
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.682 0.0 93.71 0.163 ;
      END
   END n_124393

   PIN n_124629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.786 0.0 60.814 0.163 ;
      END
   END n_124629

   PIN n_124852
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.714 0.0 89.742 0.163 ;
      END
   END n_124852

   PIN n_124877
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.73 0.0 87.758 0.163 ;
      END
   END n_124877

   PIN n_125649
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.066 0.0 78.094 0.163 ;
      END
   END n_125649

   PIN n_126016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.066 154.717 30.094 154.88 ;
      END
   END n_126016

   PIN n_127097
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.946 0.0 56.974 0.163 ;
      END
   END n_127097

   PIN n_127103
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.802 0.0 66.83 0.163 ;
      END
   END n_127103

   PIN n_127612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.586 0.0 97.614 0.163 ;
      END
   END n_127612

   PIN n_128902
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.106 154.717 37.134 154.88 ;
      END
   END n_128902

   PIN n_129209
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 64.69 0.0 64.718 0.163 ;
      END
   END n_129209

   PIN n_129975
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 91.506 0.163 91.534 ;
      END
   END n_129975

   PIN n_133431
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.394 154.717 121.422 154.88 ;
      END
   END n_133431

   PIN n_134167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.81 0.0 37.838 0.163 ;
      END
   END n_134167

   PIN n_134694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.722 0.163 60.75 ;
      END
   END n_134694

   PIN n_13477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.09 0.0 143.118 0.163 ;
      END
   END n_13477

   PIN n_13502
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 191.41 0.0 191.438 0.163 ;
      END
   END n_13502

   PIN n_137787
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 153.074 154.717 153.102 154.88 ;
      END
   END n_137787

   PIN n_137874
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.138 0.0 161.166 0.163 ;
      END
   END n_137874

   PIN n_143007
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.986 154.717 48.014 154.88 ;
      END
   END n_143007

   PIN n_144214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.314 0.0 163.342 0.163 ;
      END
   END n_144214

   PIN n_16610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.258 154.717 142.286 154.88 ;
      END
   END n_16610

   PIN n_16611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.45 154.717 142.478 154.88 ;
      END
   END n_16611

   PIN n_18394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 4.786 248.0 4.814 ;
      END
   END n_18394

   PIN n_18395
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 49.266 248.0 49.294 ;
      END
   END n_18395

   PIN n_18396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 45.298 248.0 45.326 ;
      END
   END n_18396

   PIN n_18397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 37.682 248.0 37.71 ;
      END
   END n_18397

   PIN n_18398
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 175.538 0.0 175.566 0.163 ;
      END
   END n_18398

   PIN n_18400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 170.482 0.0 170.51 0.163 ;
      END
   END n_18400

   PIN n_18779
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 45.234 248.0 45.262 ;
      END
   END n_18779

   PIN n_19896
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 234.802 0.0 234.83 0.163 ;
      END
   END n_19896

   PIN n_19897
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 4.722 248.0 4.75 ;
      END
   END n_19897

   PIN n_19898
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 193.586 0.0 193.614 0.163 ;
      END
   END n_19898

   PIN n_19899
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 193.522 0.0 193.55 0.163 ;
      END
   END n_19899

   PIN n_20359
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 14.642 248.0 14.67 ;
      END
   END n_20359

   PIN n_20449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 200.498 154.717 200.526 154.88 ;
      END
   END n_20449

   PIN n_20564
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 175.026 0.0 175.054 0.163 ;
      END
   END n_20564

   PIN n_20565
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.274 0.0 172.302 0.163 ;
      END
   END n_20565

   PIN n_20644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 183.922 0.0 183.95 0.163 ;
      END
   END n_20644

   PIN n_20800
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.034 0.0 186.062 0.163 ;
      END
   END n_20800

   PIN n_21064
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.954 154.717 147.982 154.88 ;
      END
   END n_21064

   PIN n_21065
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 175.986 154.717 176.014 154.88 ;
      END
   END n_21065

   PIN n_21066
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.762 154.717 211.79 154.88 ;
      END
   END n_21066

   PIN n_21069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 175.922 154.717 175.95 154.88 ;
      END
   END n_21069

   PIN n_21096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 63.09 248.0 63.118 ;
      END
   END n_21096

   PIN n_21097
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 56.882 248.0 56.91 ;
      END
   END n_21097

   PIN n_21145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 43.826 248.0 43.854 ;
      END
   END n_21145

   PIN n_21358
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.322 154.717 142.35 154.88 ;
      END
   END n_21358

   PIN n_21365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 56.946 248.0 56.974 ;
      END
   END n_21365

   PIN n_21400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 141.362 154.717 141.39 154.88 ;
      END
   END n_21400

   PIN n_21449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.402 154.717 164.43 154.88 ;
      END
   END n_21449

   PIN n_21451
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.322 0.0 182.35 0.163 ;
      END
   END n_21451

   PIN n_21616
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 14.322 248.0 14.35 ;
      END
   END n_21616

   PIN n_21617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 10.738 248.0 10.766 ;
      END
   END n_21617

   PIN n_21621
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 30.194 248.0 30.222 ;
      END
   END n_21621

   PIN n_21671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 244.786 0.0 244.814 0.163 ;
      END
   END n_21671

   PIN n_21890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 10.866 248.0 10.894 ;
      END
   END n_21890

   PIN n_22137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 72.69 248.0 72.718 ;
      END
   END n_22137

   PIN n_22166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 30.002 248.0 30.03 ;
      END
   END n_22166

   PIN n_22167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 33.522 248.0 33.55 ;
      END
   END n_22167

   PIN n_22235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 201.714 0.0 201.742 0.163 ;
      END
   END n_22235

   PIN n_22448
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 240.114 0.0 240.142 0.163 ;
      END
   END n_22448

   PIN n_22449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 24.242 248.0 24.27 ;
      END
   END n_22449

   PIN n_22475
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 26.162 248.0 26.19 ;
      END
   END n_22475

   PIN n_22476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 43.762 248.0 43.79 ;
      END
   END n_22476

   PIN n_22516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 237.042 0.0 237.07 0.163 ;
      END
   END n_22516

   PIN n_22541
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 30.13 248.0 30.158 ;
      END
   END n_22541

   PIN n_22817
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.146 0.0 172.174 0.163 ;
      END
   END n_22817

   PIN n_23018
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 34.354 248.0 34.382 ;
      END
   END n_23018

   PIN n_23041
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.154 0.0 143.182 0.163 ;
      END
   END n_23041

   PIN n_23125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 91.314 248.0 91.342 ;
      END
   END n_23125

   PIN n_23330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 101.362 248.0 101.39 ;
      END
   END n_23330

   PIN n_23555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.442 0.0 139.47 0.163 ;
      END
   END n_23555

   PIN n_23647
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 91.762 248.0 91.79 ;
      END
   END n_23647

   PIN n_23667
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.626 0.0 160.654 0.163 ;
      END
   END n_23667

   PIN n_23669
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.682 0.0 133.71 0.163 ;
      END
   END n_23669

   PIN n_23722
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.746 0.0 133.774 0.163 ;
      END
   END n_23722

   PIN n_23768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 87.538 248.0 87.566 ;
      END
   END n_23768

   PIN n_24318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.562 0.0 160.59 0.163 ;
      END
   END n_24318

   PIN n_24395
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 120.754 248.0 120.782 ;
      END
   END n_24395

   PIN n_24709
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.458 0.0 201.486 0.163 ;
      END
   END n_24709

   PIN n_25046
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 87.666 248.0 87.694 ;
      END
   END n_25046

   PIN n_26039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 206.962 0.0 206.99 0.163 ;
      END
   END n_26039

   PIN n_26266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 233.65 0.0 233.678 0.163 ;
      END
   END n_26266

   PIN n_26268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 225.714 0.0 225.742 0.163 ;
      END
   END n_26268

   PIN n_26406
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 99.186 248.0 99.214 ;
      END
   END n_26406

   PIN n_26895
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.834 0.0 230.862 0.163 ;
      END
   END n_26895

   PIN n_26897
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 237.426 0.0 237.454 0.163 ;
      END
   END n_26897

   PIN n_26908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 202.802 0.0 202.83 0.163 ;
      END
   END n_26908

   PIN n_27622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 191.41 154.717 191.438 154.88 ;
      END
   END n_27622

   PIN n_27970
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 192.754 0.0 192.782 0.163 ;
      END
   END n_27970

   PIN n_27972
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 187.762 0.0 187.79 0.163 ;
      END
   END n_27972

   PIN n_2799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.29 0.0 26.318 0.163 ;
      END
   END n_2799

   PIN n_28572
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 145.33 248.0 145.358 ;
      END
   END n_28572

   PIN n_28574
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 145.266 248.0 145.294 ;
      END
   END n_28574

   PIN n_2861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 175.154 154.717 175.182 154.88 ;
      END
   END n_2861

   PIN n_2871
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.61 0.0 138.638 0.163 ;
      END
   END n_2871

   PIN n_28733
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 150.002 248.0 150.03 ;
      END
   END n_28733

   PIN n_29056
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.57 154.717 227.598 154.88 ;
      END
   END n_29056

   PIN n_29058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.378 154.717 227.406 154.88 ;
      END
   END n_29058

   PIN n_32114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.306 154.717 80.334 154.88 ;
      END
   END n_32114

   PIN n_32115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.114 154.717 80.142 154.88 ;
      END
   END n_32115

   PIN n_32440
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.762 154.717 83.79 154.88 ;
      END
   END n_32440

   PIN n_32718
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.258 154.717 38.286 154.88 ;
      END
   END n_32718

   PIN n_32740
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.378 154.717 51.406 154.88 ;
      END
   END n_32740

   PIN n_32741
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.186 154.717 51.214 154.88 ;
      END
   END n_32741

   PIN n_32769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.618 154.717 69.646 154.88 ;
      END
   END n_32769

   PIN n_33082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.682 154.717 61.71 154.88 ;
      END
   END n_33082

   PIN n_33167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.954 154.717 43.982 154.88 ;
      END
   END n_33167

   PIN n_33364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.89 154.717 75.918 154.88 ;
      END
   END n_33364

   PIN n_33881
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.602 154.717 87.63 154.88 ;
      END
   END n_33881

   PIN n_34014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.506 154.717 3.534 154.88 ;
      END
   END n_34014

   PIN n_34377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.586 154.717 41.614 154.88 ;
      END
   END n_34377

   PIN n_34609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 80.242 154.717 80.27 154.88 ;
      END
   END n_34609

   PIN n_34610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.434 154.717 80.462 154.88 ;
      END
   END n_34610

   PIN n_34731
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 87.666 154.717 87.694 154.88 ;
      END
   END n_34731

   PIN n_34808
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.522 154.717 41.55 154.88 ;
      END
   END n_34808

   PIN n_3513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.21 154.717 172.238 154.88 ;
      END
   END n_3513

   PIN n_35434
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.77 154.717 54.798 154.88 ;
      END
   END n_35434

   PIN n_36613
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.626 154.717 64.654 154.88 ;
      END
   END n_36613

   PIN n_37477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.33 154.717 25.358 154.88 ;
      END
   END n_37477

   PIN n_37556
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.314 154.717 91.342 154.88 ;
      END
   END n_37556

   PIN n_37622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.73 154.717 87.758 154.88 ;
      END
   END n_37622

   PIN n_37665
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.346 154.717 95.374 154.88 ;
      END
   END n_37665

   PIN n_37690
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.858 154.717 79.886 154.88 ;
      END
   END n_37690

   PIN n_382
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.818 154.717 152.846 154.88 ;
      END
   END n_382

   PIN n_39240
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.978 154.717 69.006 154.88 ;
      END
   END n_39240

   PIN n_39453
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.09 0.0 103.118 0.163 ;
      END
   END n_39453

   PIN n_39845
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.93 154.717 106.958 154.88 ;
      END
   END n_39845

   PIN n_40155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.918 24.114 248.0 24.142 ;
      END
   END n_40155

   PIN n_40158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 82.162 248.0 82.19 ;
      END
   END n_40158

   PIN n_40330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 53.362 248.0 53.39 ;
      END
   END n_40330

   PIN n_40445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 240.242 0.0 240.27 0.163 ;
      END
   END n_40445

   PIN n_40476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 246.834 0.0 246.862 0.163 ;
      END
   END n_40476

   PIN n_40561
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 223.986 0.0 224.014 0.163 ;
      END
   END n_40561

   PIN n_40564
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.442 0.0 235.47 0.163 ;
      END
   END n_40564

   PIN n_40626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 223.922 0.0 223.95 0.163 ;
      END
   END n_40626

   PIN n_40648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 241.394 0.0 241.422 0.163 ;
      END
   END n_40648

   PIN n_40695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 210.61 0.0 210.638 0.163 ;
      END
   END n_40695

   PIN n_40706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 72.626 248.0 72.654 ;
      END
   END n_40706

   PIN n_40727
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 222.386 0.0 222.414 0.163 ;
      END
   END n_40727

   PIN n_48178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.034 154.717 74.062 154.88 ;
      END
   END n_48178

   PIN n_48510
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.242 154.717 16.27 154.88 ;
      END
   END n_48510

   PIN n_48907
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.426 154.717 77.454 154.88 ;
      END
   END n_48907

   PIN n_49236
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.722 0.0 228.75 0.163 ;
      END
   END n_49236

   PIN n_5058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.578 0.0 150.606 0.163 ;
      END
   END n_5058

   PIN n_5059
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.77 0.0 150.798 0.163 ;
      END
   END n_5059

   PIN n_5115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.17 154.717 149.198 154.88 ;
      END
   END n_5115

   PIN n_51768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.114 154.717 72.142 154.88 ;
      END
   END n_51768

   PIN n_54235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.362 154.717 77.39 154.88 ;
      END
   END n_54235

   PIN n_54706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 63.026 248.0 63.054 ;
      END
   END n_54706

   PIN n_5505
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.746 154.717 133.774 154.88 ;
      END
   END n_5505

   PIN n_5571
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.93 0.0 162.958 0.163 ;
      END
   END n_5571

   PIN n_57100
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.234 154.717 77.262 154.88 ;
      END
   END n_57100

   PIN n_58492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 247.837 62.962 248.0 62.99 ;
      END
   END n_58492

   PIN n_58941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.37 154.717 72.398 154.88 ;
      END
   END n_58941

   PIN n_60391
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.698 0.0 235.726 0.163 ;
      END
   END n_60391

   PIN n_6364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.146 154.717 172.174 154.88 ;
      END
   END n_6364

   PIN n_63870
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 219.506 0.0 219.534 0.163 ;
      END
   END n_63870

   PIN n_6635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.946 154.717 152.974 154.88 ;
      END
   END n_6635

   PIN n_7003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.898 0.0 246.926 0.163 ;
      END
   END n_7003

   PIN n_7337
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 172.21 154.717 172.238 154.88 ;
      END
   END n_7337

   PIN n_7696
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.85 0.163 60.878 ;
      END
   END n_7696

   PIN n_7848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.194 154.717 166.222 154.88 ;
      END
   END n_7848

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 248.0 154.88 ;
      LAYER V1 ;
         RECT 0.0 0.0 248.0 154.88 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 248.0 154.88 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 248.0 154.88 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 248.0 154.88 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 248.0 154.88 ;
      LAYER M1 ;
         RECT 0.0 0.0 248.0 154.88 ;
   END
END h1_mgc_matrix_mult_a

MACRO h0_mgc_matrix_mult_a
   CLASS BLOCK ;
   FOREIGN h0 ;
   ORIGIN 0 0 ;
   SIZE 241.856 BY 122.24 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN10233_b_2_6_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.218 122.077 135.246 122.24 ;
      END
   END FE_OFN10233_b_2_6_0

   PIN FE_OFN10257_b_2_4_6
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.578 122.077 150.606 122.24 ;
      END
   END FE_OFN10257_b_2_4_6

   PIN FE_OFN10260_b_2_4_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.946 122.077 128.974 122.24 ;
      END
   END FE_OFN10260_b_2_4_5

   PIN FE_OFN10293_b_2_2_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.306 122.077 88.334 122.24 ;
      END
   END FE_OFN10293_b_2_2_3

   PIN FE_OFN1071_n_16034
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 98.546 241.856 98.574 ;
      END
   END FE_OFN1071_n_16034

   PIN FE_OFN1086_n_21187
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.962 122.077 230.99 122.24 ;
      END
   END FE_OFN1086_n_21187

   PIN FE_OFN11430_n_142905
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 106.226 241.856 106.254 ;
      END
   END FE_OFN11430_n_142905

   PIN FE_OFN11434_n_142919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 109.81 241.856 109.838 ;
      END
   END FE_OFN11434_n_142919

   PIN FE_OFN11435_n_142919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.434 122.077 112.462 122.24 ;
      END
   END FE_OFN11435_n_142919

   PIN FE_OFN1157_n_10648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.858 122.077 207.886 122.24 ;
      END
   END FE_OFN1157_n_10648

   PIN FE_OFN11706_n_142947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 177.714 122.077 177.742 122.24 ;
      END
   END FE_OFN11706_n_142947

   PIN FE_OFN11707_n_142947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 110.066 241.856 110.094 ;
      END
   END FE_OFN11707_n_142947

   PIN FE_OFN12301_n_111727
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 102.898 241.856 102.926 ;
      END
   END FE_OFN12301_n_111727

   PIN FE_OFN12386_n_142906
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.706 122.077 150.734 122.24 ;
      END
   END FE_OFN12386_n_142906

   PIN FE_OFN12400_n_694
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.594 122.077 100.622 122.24 ;
      END
   END FE_OFN12400_n_694

   PIN FE_OFN12617_n_112689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.002 122.077 134.03 122.24 ;
      END
   END FE_OFN12617_n_112689

   PIN FE_OFN12618_n_112689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 146.802 122.077 146.83 122.24 ;
      END
   END FE_OFN12618_n_112689

   PIN FE_OFN13018_n_142950
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.706 122.077 158.734 122.24 ;
      END
   END FE_OFN13018_n_142950

   PIN FE_OFN15062_n_12711
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.25 122.077 131.278 122.24 ;
      END
   END FE_OFN15062_n_12711

   PIN FE_OFN15077_n_14458
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.146 122.077 180.174 122.24 ;
      END
   END FE_OFN15077_n_14458

   PIN FE_OFN15252_n_39084
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 223.73 122.077 223.758 122.24 ;
      END
   END FE_OFN15252_n_39084

   PIN FE_OFN15923_n_143045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 115.058 241.856 115.086 ;
      END
   END FE_OFN15923_n_143045

   PIN FE_OFN15925_n_112550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.186 122.077 139.214 122.24 ;
      END
   END FE_OFN15925_n_112550

   PIN FE_OFN15930_n_143241
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.178 122.077 112.206 122.24 ;
      END
   END FE_OFN15930_n_143241

   PIN FE_OFN16294_delay_add_ln34_unr2_unr3_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.858 122.077 159.886 122.24 ;
      END
   END FE_OFN16294_delay_add_ln34_unr2_unr3_stage2_stallmux_q_15_

   PIN FE_OFN16366_b_2_4_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.778 122.077 169.806 122.24 ;
      END
   END FE_OFN16366_b_2_4_1

   PIN FE_OFN16771_n_16098
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 118.194 241.856 118.222 ;
      END
   END FE_OFN16771_n_16098

   PIN FE_OFN17162_n_132699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.45 122.077 62.478 122.24 ;
      END
   END FE_OFN17162_n_132699

   PIN FE_OFN17165_n_134675
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.29 122.077 162.318 122.24 ;
      END
   END FE_OFN17165_n_134675

   PIN FE_OFN17200_n_16166
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.402 122.077 196.43 122.24 ;
      END
   END FE_OFN17200_n_16166

   PIN FE_OFN17265_n_140245
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 114.098 241.856 114.126 ;
      END
   END FE_OFN17265_n_140245

   PIN FE_OFN18609_b_2_2_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.858 122.077 111.886 122.24 ;
      END
   END FE_OFN18609_b_2_2_0

   PIN FE_OFN18810_n_143645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.554 122.077 181.582 122.24 ;
      END
   END FE_OFN18810_n_143645

   PIN FE_OFN19059_n_19681
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.698 122.077 227.726 122.24 ;
      END
   END FE_OFN19059_n_19681

   PIN FE_OFN19145_n_143045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 110.578 241.856 110.606 ;
      END
   END FE_OFN19145_n_143045

   PIN FE_OFN19307_b_2_2_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.026 122.077 135.054 122.24 ;
      END
   END FE_OFN19307_b_2_2_1

   PIN FE_OFN2160_n_19626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.298 122.077 229.326 122.24 ;
      END
   END FE_OFN2160_n_19626

   PIN FE_OFN2283_n_19629
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.322 122.077 158.35 122.24 ;
      END
   END FE_OFN2283_n_19629

   PIN FE_OFN3286_n_117368
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.802 122.077 146.83 122.24 ;
      END
   END FE_OFN3286_n_117368

   PIN FE_OFN3294_n_8246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 94.578 241.856 94.606 ;
      END
   END FE_OFN3294_n_8246

   PIN FE_OFN3442_n_12341
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 117.938 241.856 117.966 ;
      END
   END FE_OFN3442_n_12341

   PIN FE_OFN3574_n_133235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.234 122.077 85.262 122.24 ;
      END
   END FE_OFN3574_n_133235

   PIN FE_OFN3613_n_112427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.698 122.077 115.726 122.24 ;
      END
   END FE_OFN3613_n_112427

   PIN FE_OFN3656_n_112550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.314 122.077 123.342 122.24 ;
      END
   END FE_OFN3656_n_112550

   PIN FE_OFN3723_n_143241
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.922 122.077 111.95 122.24 ;
      END
   END FE_OFN3723_n_143241

   PIN FE_OFN606_n_8387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 240.818 122.077 240.846 122.24 ;
      END
   END FE_OFN606_n_8387

   PIN FE_OFN703_n_21657
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.346 122.077 231.374 122.24 ;
      END
   END FE_OFN703_n_21657

   PIN FE_OFN757_n_21703
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.658 122.077 204.686 122.24 ;
      END
   END FE_OFN757_n_21703

   PIN FE_OFN797_n_21129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.09 122.077 239.118 122.24 ;
      END
   END FE_OFN797_n_21129

   PIN add_5900_51_n_148
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 55.218 241.856 55.246 ;
      END
   END add_5900_51_n_148

   PIN add_5900_51_n_77
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.722 122.077 172.75 122.24 ;
      END
   END add_5900_51_n_77

   PIN delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 166.642 122.077 166.67 122.24 ;
      END
   END delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_

   PIN delay_add_ln34_unr2_unr2_stage2_stallmux_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 193.01 122.077 193.038 122.24 ;
      END
   END delay_add_ln34_unr2_unr2_stage2_stallmux_z_12_

   PIN delay_add_ln34_unr2_unr3_stage2_stallmux_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 199.986 122.077 200.014 122.24 ;
      END
   END delay_add_ln34_unr2_unr3_stage2_stallmux_q_10_

   PIN delay_add_ln34_unr2_unr3_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 102.834 241.856 102.862 ;
      END
   END delay_add_ln34_unr2_unr3_stage2_stallmux_q_3_

   PIN delay_add_ln34_unr2_unr3_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 118.258 241.856 118.286 ;
      END
   END delay_add_ln34_unr2_unr3_stage2_stallmux_q_4_

   PIN delay_add_ln34_unr2_unr3_stage2_stallmux_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 113.842 241.856 113.87 ;
      END
   END delay_add_ln34_unr2_unr3_stage2_stallmux_q_8_

   PIN delay_add_ln34_unr2_unr5_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 212.274 122.077 212.302 122.24 ;
      END
   END delay_add_ln34_unr2_unr5_stage2_stallmux_q_14_

   PIN delay_add_ln34_unr2_unr5_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 105.97 241.856 105.998 ;
      END
   END delay_add_ln34_unr2_unr5_stage2_stallmux_q_7_

   PIN delay_add_ln34_unr2_unr5_stage2_stallmux_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 109.874 241.856 109.902 ;
      END
   END delay_add_ln34_unr2_unr5_stage2_stallmux_q_8_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.778 122.077 201.806 122.24 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_3_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 189.106 122.077 189.134 122.24 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_4_

   PIN delay_add_ln34_unr2_unr8_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 90.674 241.856 90.702 ;
      END
   END delay_add_ln34_unr2_unr8_stage2_stallmux_q_3_

   PIN mul_4665_72_n_202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.162 122.077 66.19 122.24 ;
      END
   END mul_4665_72_n_202

   PIN mul_4665_72_n_221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.722 122.077 20.75 122.24 ;
      END
   END mul_4665_72_n_221

   PIN mul_4665_72_n_230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.626 122.077 104.654 122.24 ;
      END
   END mul_4665_72_n_230

   PIN mul_4665_72_n_295
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.402 122.077 4.43 122.24 ;
      END
   END mul_4665_72_n_295

   PIN mul_4665_72_n_337
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.346 122.077 39.374 122.24 ;
      END
   END mul_4665_72_n_337

   PIN mul_4665_72_n_848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.066 122.077 70.094 122.24 ;
      END
   END mul_4665_72_n_848

   PIN mul_4667_72_n_184
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 181.49 122.077 181.518 122.24 ;
      END
   END mul_4667_72_n_184

   PIN mul_4667_72_n_265
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 185.33 122.077 185.358 122.24 ;
      END
   END mul_4667_72_n_265

   PIN mul_4667_72_n_304
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.778 122.077 113.806 122.24 ;
      END
   END mul_4667_72_n_304

   PIN mul_4667_72_n_308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.37 122.077 128.398 122.24 ;
      END
   END mul_4667_72_n_308

   PIN mul_4667_72_n_316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.65 122.077 81.678 122.24 ;
      END
   END mul_4667_72_n_316

   PIN mul_4667_72_n_323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.45 122.077 78.478 122.24 ;
      END
   END mul_4667_72_n_323

   PIN mul_4667_72_n_324
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.682 122.077 77.71 122.24 ;
      END
   END mul_4667_72_n_324

   PIN mul_4667_72_n_327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.81 122.077 77.838 122.24 ;
      END
   END mul_4667_72_n_327

   PIN mul_4667_72_n_66
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 158.45 122.077 158.478 122.24 ;
      END
   END mul_4667_72_n_66

   PIN mul_4669_72_n_225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 135.282 122.077 135.31 122.24 ;
      END
   END mul_4669_72_n_225

   PIN mul_4669_72_n_304
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.978 122.077 125.006 122.24 ;
      END
   END mul_4669_72_n_304

   PIN mul_4669_72_n_314
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.834 122.077 118.862 122.24 ;
      END
   END mul_4669_72_n_314

   PIN mul_4669_72_n_316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.906 122.077 121.934 122.24 ;
      END
   END mul_4669_72_n_316

   PIN mul_4669_72_n_66
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 185.33 122.077 185.358 122.24 ;
      END
   END mul_4669_72_n_66

   PIN mul_ln34_unr0_unr6_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.482 241.856 90.51 ;
      END
   END mul_ln34_unr0_unr6_z_14_

   PIN mul_ln34_unr2_unr2_z_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 106.034 241.856 106.062 ;
      END
   END mul_ln34_unr2_unr2_z_0_

   PIN mul_ln34_unr2_unr2_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 63.73 241.856 63.758 ;
      END
   END mul_ln34_unr2_unr2_z_14_

   PIN mul_ln34_unr2_unr2_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.154 122.077 239.182 122.24 ;
      END
   END mul_ln34_unr2_unr2_z_7_

   PIN n_10378
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.866 122.077 146.894 122.24 ;
      END
   END n_10378

   PIN n_10669
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.946 122.077 120.974 122.24 ;
      END
   END n_10669

   PIN n_11011
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 86.77 241.856 86.798 ;
      END
   END n_11011

   PIN n_111968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 223.666 122.077 223.694 122.24 ;
      END
   END n_111968

   PIN n_112778
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 55.922 241.856 55.95 ;
      END
   END n_112778

   PIN n_112779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 55.986 241.856 56.014 ;
      END
   END n_112779

   PIN n_112812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 52.082 241.856 52.11 ;
      END
   END n_112812

   PIN n_112817
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.338 122.077 164.366 122.24 ;
      END
   END n_112817

   PIN n_112831
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 53.49 241.856 53.518 ;
      END
   END n_112831

   PIN n_112845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 46.258 241.856 46.286 ;
      END
   END n_112845

   PIN n_112880
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 46.258 241.856 46.286 ;
      END
   END n_112880

   PIN n_112890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.586 122.077 81.614 122.24 ;
      END
   END n_112890

   PIN n_112959
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.778 122.077 73.806 122.24 ;
      END
   END n_112959

   PIN n_113054
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.314 241.856 75.342 ;
      END
   END n_113054

   PIN n_113100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.498 122.077 72.526 122.24 ;
      END
   END n_113100

   PIN n_113160
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.882 122.077 96.91 122.24 ;
      END
   END n_113160

   PIN n_113191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.97 122.077 169.998 122.24 ;
      END
   END n_113191

   PIN n_113195
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 56.05 241.856 56.078 ;
      END
   END n_113195

   PIN n_113217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 32.818 241.856 32.846 ;
      END
   END n_113217

   PIN n_113223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.746 122.077 149.774 122.24 ;
      END
   END n_113223

   PIN n_113308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.09 122.077 143.118 122.24 ;
      END
   END n_113308

   PIN n_113317
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.73 122.077 143.758 122.24 ;
      END
   END n_113317

   PIN n_113342
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.906 122.077 89.934 122.24 ;
      END
   END n_113342

   PIN n_113343
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.778 122.077 89.806 122.24 ;
      END
   END n_113343

   PIN n_113447
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 173.81 122.077 173.838 122.24 ;
      END
   END n_113447

   PIN n_113479
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 25.458 241.856 25.486 ;
      END
   END n_113479

   PIN n_113480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.842 122.077 97.87 122.24 ;
      END
   END n_113480

   PIN n_113481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.914 122.077 92.942 122.24 ;
      END
   END n_113481

   PIN n_113503
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.234 122.077 93.262 122.24 ;
      END
   END n_113503

   PIN n_113516
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.842 122.077 89.87 122.24 ;
      END
   END n_113516

   PIN n_113517
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.714 122.077 89.742 122.24 ;
      END
   END n_113517

   PIN n_113545
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.53 122.077 172.558 122.24 ;
      END
   END n_113545

   PIN n_113830
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 17.97 241.856 17.998 ;
      END
   END n_113830

   PIN n_113933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.954 122.077 155.982 122.24 ;
      END
   END n_113933

   PIN n_113934
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.77 122.077 150.798 122.24 ;
      END
   END n_113934

   PIN n_114134
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.658 122.077 100.686 122.24 ;
      END
   END n_114134

   PIN n_114136
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.002 122.077 70.03 122.24 ;
      END
   END n_114136

   PIN n_114331
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.042 122.077 125.07 122.24 ;
      END
   END n_114331

   PIN n_114597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 153.458 122.077 153.486 122.24 ;
      END
   END n_114597

   PIN n_114598
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.834 122.077 150.862 122.24 ;
      END
   END n_114598

   PIN n_114821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.842 122.077 113.87 122.24 ;
      END
   END n_114821

   PIN n_114951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.658 122.077 116.686 122.24 ;
      END
   END n_114951

   PIN n_115117
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.794 122.077 71.822 122.24 ;
      END
   END n_115117

   PIN n_115119
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.954 122.077 91.982 122.24 ;
      END
   END n_115119

   PIN n_115219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.826 122.077 123.854 122.24 ;
      END
   END n_115219

   PIN n_116269
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.426 122.077 85.454 122.24 ;
      END
   END n_116269

   PIN n_116470
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.306 122.077 112.334 122.24 ;
      END
   END n_116470

   PIN n_117525
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 48.242 241.856 48.27 ;
      END
   END n_117525

   PIN n_117559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 29.618 241.856 29.646 ;
      END
   END n_117559

   PIN n_117560
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 32.242 241.856 32.27 ;
      END
   END n_117560

   PIN n_117582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.842 122.077 73.87 122.24 ;
      END
   END n_117582

   PIN n_117603
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.138 122.077 81.166 122.24 ;
      END
   END n_117603

   PIN n_117620
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.994 122.077 147.022 122.24 ;
      END
   END n_117620

   PIN n_118017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.842 122.077 57.87 122.24 ;
      END
   END n_118017

   PIN n_118035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.522 241.856 25.55 ;
      END
   END n_118035

   PIN n_118166
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.146 122.077 84.174 122.24 ;
      END
   END n_118166

   PIN n_118364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.394 122.077 153.422 122.24 ;
      END
   END n_118364

   PIN n_119552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.682 122.077 117.71 122.24 ;
      END
   END n_119552

   PIN n_119619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 40.754 241.856 40.782 ;
      END
   END n_119619

   PIN n_119690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.418 122.077 66.446 122.24 ;
      END
   END n_119690

   PIN n_119691
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.122 122.077 67.15 122.24 ;
      END
   END n_119691

   PIN n_119709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.514 122.077 62.542 122.24 ;
      END
   END n_119709

   PIN n_119812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.01 122.077 97.038 122.24 ;
      END
   END n_119812

   PIN n_119886
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 20.978 241.856 21.006 ;
      END
   END n_119886

   PIN n_119969
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.282 122.077 159.31 122.24 ;
      END
   END n_119969

   PIN n_120042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.458 122.077 169.486 122.24 ;
      END
   END n_120042

   PIN n_120044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.57 122.077 51.598 122.24 ;
      END
   END n_120044

   PIN n_120045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.562 122.077 56.59 122.24 ;
      END
   END n_120045

   PIN n_120129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.914 122.077 100.942 122.24 ;
      END
   END n_120129

   PIN n_120131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.266 122.077 89.294 122.24 ;
      END
   END n_120131

   PIN n_120499
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.61 122.077 58.638 122.24 ;
      END
   END n_120499

   PIN n_120794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.786 122.077 36.814 122.24 ;
      END
   END n_120794

   PIN n_121083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.474 122.077 31.502 122.24 ;
      END
   END n_121083

   PIN n_121084
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.378 122.077 35.406 122.24 ;
      END
   END n_121084

   PIN n_121196
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.866 241.856 90.894 ;
      END
   END n_121196

   PIN n_121291
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 85.362 241.856 85.39 ;
      END
   END n_121291

   PIN n_121522
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 94.642 241.856 94.67 ;
      END
   END n_121522

   PIN n_121732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 37.298 241.856 37.326 ;
      END
   END n_121732

   PIN n_121779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.026 122.077 63.054 122.24 ;
      END
   END n_121779

   PIN n_121908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.05 122.077 8.078 122.24 ;
      END
   END n_121908

   PIN n_121917
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.594 122.077 132.622 122.24 ;
      END
   END n_121917

   PIN n_121918
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.474 122.077 135.502 122.24 ;
      END
   END n_121918

   PIN n_122005
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.042 122.077 101.07 122.24 ;
      END
   END n_122005

   PIN n_122026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.506 122.077 147.534 122.24 ;
      END
   END n_122026

   PIN n_122106
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.666 122.077 31.694 122.24 ;
      END
   END n_122106

   PIN n_122300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.282 122.077 79.31 122.24 ;
      END
   END n_122300

   PIN n_122476
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.378 241.856 75.406 ;
      END
   END n_122476

   PIN n_122532
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 53.746 241.856 53.774 ;
      END
   END n_122532

   PIN n_123300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.058 122.077 91.086 122.24 ;
      END
   END n_123300

   PIN n_123316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.434 122.077 120.462 122.24 ;
      END
   END n_123316

   PIN n_123618
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.762 122.077 75.79 122.24 ;
      END
   END n_123618

   PIN n_123955
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 56.114 241.856 56.142 ;
      END
   END n_123955

   PIN n_124058
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.914 122.077 100.942 122.24 ;
      END
   END n_124058

   PIN n_124589
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.594 122.077 60.622 122.24 ;
      END
   END n_124589

   PIN n_124590
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.578 122.077 62.606 122.24 ;
      END
   END n_124590

   PIN n_124859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 86.834 241.856 86.862 ;
      END
   END n_124859

   PIN n_125049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 60.146 241.856 60.174 ;
      END
   END n_125049

   PIN n_125190
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 83.186 241.856 83.214 ;
      END
   END n_125190

   PIN n_125260
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 82.866 241.856 82.894 ;
      END
   END n_125260

   PIN n_125261
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 82.738 241.856 82.766 ;
      END
   END n_125261

   PIN n_125371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.73 122.077 31.758 122.24 ;
      END
   END n_125371

   PIN n_125378
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.73 122.077 127.758 122.24 ;
      END
   END n_125378

   PIN n_125536
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 85.938 241.856 85.966 ;
      END
   END n_125536

   PIN n_125537
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 83.442 241.856 83.47 ;
      END
   END n_125537

   PIN n_125551
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 143.09 122.077 143.118 122.24 ;
      END
   END n_125551

   PIN n_12570
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.114 122.077 152.142 122.24 ;
      END
   END n_12570

   PIN n_125714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 78.962 241.856 78.99 ;
      END
   END n_125714

   PIN n_125785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 73.202 122.077 73.23 122.24 ;
      END
   END n_125785

   PIN n_126191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.682 122.077 77.71 122.24 ;
      END
   END n_126191

   PIN n_126306
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 69.234 241.856 69.262 ;
      END
   END n_126306

   PIN n_126307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 69.298 241.856 69.326 ;
      END
   END n_126307

   PIN n_126587
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.722 122.077 60.75 122.24 ;
      END
   END n_126587

   PIN n_126600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.506 122.077 75.534 122.24 ;
      END
   END n_126600

   PIN n_126601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.642 122.077 70.67 122.24 ;
      END
   END n_126601

   PIN n_12712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.186 122.077 131.214 122.24 ;
      END
   END n_12712

   PIN n_127297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.562 122.077 64.59 122.24 ;
      END
   END n_127297

   PIN n_127737
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 67.698 241.856 67.726 ;
      END
   END n_127737

   PIN n_127742
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.442 241.856 75.47 ;
      END
   END n_127742

   PIN n_127891
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.626 122.077 48.654 122.24 ;
      END
   END n_127891

   PIN n_128372
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.402 122.077 60.43 122.24 ;
      END
   END n_128372

   PIN n_128584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 62.258 241.856 62.286 ;
      END
   END n_128584

   PIN n_128848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 77.618 241.856 77.646 ;
      END
   END n_128848

   PIN n_128849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.506 241.856 75.534 ;
      END
   END n_128849

   PIN n_128989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.058 122.077 75.086 122.24 ;
      END
   END n_128989

   PIN n_129129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 146.866 122.077 146.894 122.24 ;
      END
   END n_129129

   PIN n_129403
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.13 122.077 62.158 122.24 ;
      END
   END n_129403

   PIN n_129491
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 4.914 241.856 4.942 ;
      END
   END n_129491

   PIN n_129545
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.002 122.077 38.03 122.24 ;
      END
   END n_129545

   PIN n_129619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 62.258 241.856 62.286 ;
      END
   END n_129619

   PIN n_129824
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.418 122.077 58.446 122.24 ;
      END
   END n_129824

   PIN n_129826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.802 122.077 50.83 122.24 ;
      END
   END n_129826

   PIN n_129827
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 4.978 241.856 5.006 ;
      END
   END n_129827

   PIN n_129828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 73.842 122.077 73.87 122.24 ;
      END
   END n_129828

   PIN n_129897
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.57 122.077 19.598 122.24 ;
      END
   END n_129897

   PIN n_130137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 40.882 241.856 40.91 ;
      END
   END n_130137

   PIN n_130202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.33 241.856 25.358 ;
      END
   END n_130202

   PIN n_130204
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.65 241.856 25.678 ;
      END
   END n_130204

   PIN n_130594
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 82.802 241.856 82.83 ;
      END
   END n_130594

   PIN n_130626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 10.098 241.856 10.126 ;
      END
   END n_130626

   PIN n_131059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 17.65 241.856 17.678 ;
      END
   END n_131059

   PIN n_131060
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 21.234 241.856 21.262 ;
      END
   END n_131060

   PIN n_131305
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.498 122.077 112.526 122.24 ;
      END
   END n_131305

   PIN n_131421
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 17.714 241.856 17.742 ;
      END
   END n_131421

   PIN n_131475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.93 122.077 146.958 122.24 ;
      END
   END n_131475

   PIN n_132026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.41 122.077 103.438 122.24 ;
      END
   END n_132026

   PIN n_132027
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.466 122.077 108.494 122.24 ;
      END
   END n_132027

   PIN n_132085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 60.978 241.856 61.006 ;
      END
   END n_132085

   PIN n_132293
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.242 122.077 112.27 122.24 ;
      END
   END n_132293

   PIN n_132825
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.786 122.077 100.814 122.24 ;
      END
   END n_132825

   PIN n_132870
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 33.138 241.856 33.166 ;
      END
   END n_132870

   PIN n_133002
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.618 122.077 109.646 122.24 ;
      END
   END n_133002

   PIN n_133183
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.162 122.077 66.19 122.24 ;
      END
   END n_133183

   PIN n_133738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.706 122.077 142.734 122.24 ;
      END
   END n_133738

   PIN n_133859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 33.01 241.856 33.038 ;
      END
   END n_133859

   PIN n_133940
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 21.426 241.856 21.454 ;
      END
   END n_133940

   PIN n_134182
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.69 122.077 104.718 122.24 ;
      END
   END n_134182

   PIN n_134553
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 33.33 241.856 33.358 ;
      END
   END n_134553

   PIN n_134648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 21.49 241.856 21.518 ;
      END
   END n_134648

   PIN n_134804
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.922 122.077 103.95 122.24 ;
      END
   END n_134804

   PIN n_135056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.018 122.077 124.046 122.24 ;
      END
   END n_135056

   PIN n_135073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.746 122.077 85.774 122.24 ;
      END
   END n_135073

   PIN n_135074
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.49 122.077 85.518 122.24 ;
      END
   END n_135074

   PIN n_135796
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 21.106 241.856 21.134 ;
      END
   END n_135796

   PIN n_135808
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 165.746 122.077 165.774 122.24 ;
      END
   END n_135808

   PIN n_136154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 10.29 241.856 10.318 ;
      END
   END n_136154

   PIN n_136201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.714 122.077 49.742 122.24 ;
      END
   END n_136201

   PIN n_136203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.914 122.077 52.942 122.24 ;
      END
   END n_136203

   PIN n_136211
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.658 122.077 52.686 122.24 ;
      END
   END n_136211

   PIN n_136212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.986 122.077 56.014 122.24 ;
      END
   END n_136212

   PIN n_136268
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 48.306 241.856 48.334 ;
      END
   END n_136268

   PIN n_136598
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 44.53 241.856 44.558 ;
      END
   END n_136598

   PIN n_136630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 48.37 241.856 48.398 ;
      END
   END n_136630

   PIN n_136660
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 71.474 241.856 71.502 ;
      END
   END n_136660

   PIN n_136842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.122 241.856 75.15 ;
      END
   END n_136842

   PIN n_136875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.298 122.077 181.326 122.24 ;
      END
   END n_136875

   PIN n_136876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 185.266 122.077 185.294 122.24 ;
      END
   END n_136876

   PIN n_136887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 178.994 122.077 179.022 122.24 ;
      END
   END n_136887

   PIN n_137597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 69.362 241.856 69.39 ;
      END
   END n_137597

   PIN n_14162
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.754 122.077 120.782 122.24 ;
      END
   END n_14162

   PIN n_143063
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.426 122.077 181.454 122.24 ;
      END
   END n_143063

   PIN n_143692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 56.882 241.856 56.91 ;
      END
   END n_143692

   PIN n_143725
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.25 122.077 139.278 122.24 ;
      END
   END n_143725

   PIN n_143810
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 71.538 241.856 71.566 ;
      END
   END n_143810

   PIN n_143811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 71.41 241.856 71.438 ;
      END
   END n_143811

   PIN n_14682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.514 122.077 118.542 122.24 ;
      END
   END n_14682

   PIN n_16033
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 94.322 241.856 94.35 ;
      END
   END n_16033

   PIN n_16164
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 59.698 241.856 59.726 ;
      END
   END n_16164

   PIN n_16207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.178 122.077 208.206 122.24 ;
      END
   END n_16207

   PIN n_16296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.922 122.077 215.95 122.24 ;
      END
   END n_16296

   PIN n_18629
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.314 122.077 235.342 122.24 ;
      END
   END n_18629

   PIN n_18630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 232.69 122.077 232.718 122.24 ;
      END
   END n_18630

   PIN n_18732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 217.074 122.077 217.102 122.24 ;
      END
   END n_18732

   PIN n_18908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.338 122.077 204.366 122.24 ;
      END
   END n_18908

   PIN n_18997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 48.434 241.856 48.462 ;
      END
   END n_18997

   PIN n_19022
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.25 122.077 235.278 122.24 ;
      END
   END n_19022

   PIN n_19642
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.026 122.077 143.054 122.24 ;
      END
   END n_19642

   PIN n_20025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 83.25 241.856 83.278 ;
      END
   END n_20025

   PIN n_20054
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 239.09 122.077 239.118 122.24 ;
      END
   END n_20054

   PIN n_20260
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 200.626 122.077 200.654 122.24 ;
      END
   END n_20260

   PIN n_20282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 154.61 122.077 154.638 122.24 ;
      END
   END n_20282

   PIN n_20329
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 40.626 241.856 40.654 ;
      END
   END n_20329

   PIN n_20334
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 173.746 122.077 173.774 122.24 ;
      END
   END n_20334

   PIN n_20442
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.402 122.077 204.43 122.24 ;
      END
   END n_20442

   PIN n_20443
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.466 122.077 204.494 122.24 ;
      END
   END n_20443

   PIN n_20690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.53 122.077 204.558 122.24 ;
      END
   END n_20690

   PIN n_20855
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 71.474 241.856 71.502 ;
      END
   END n_20855

   PIN n_20865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 67.57 241.856 67.598 ;
      END
   END n_20865

   PIN n_20867
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.594 122.077 204.622 122.24 ;
      END
   END n_20867

   PIN n_20880
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 177.522 122.077 177.55 122.24 ;
      END
   END n_20880

   PIN n_21104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 94.45 241.856 94.478 ;
      END
   END n_21104

   PIN n_21252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 56.242 241.856 56.27 ;
      END
   END n_21252

   PIN n_21408
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 231.858 122.077 231.886 122.24 ;
      END
   END n_21408

   PIN n_21512
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.082 122.077 60.11 122.24 ;
      END
   END n_21512

   PIN n_21514
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.322 122.077 62.35 122.24 ;
      END
   END n_21514

   PIN n_21917
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 98.418 241.856 98.446 ;
      END
   END n_21917

   PIN n_22013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.21 122.077 212.238 122.24 ;
      END
   END n_22013

   PIN n_22014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.914 122.077 220.942 122.24 ;
      END
   END n_22014

   PIN n_22238
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.298 122.077 85.326 122.24 ;
      END
   END n_22238

   PIN n_22308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.242 122.077 208.27 122.24 ;
      END
   END n_22308

   PIN n_22322
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.434 122.077 208.462 122.24 ;
      END
   END n_22322

   PIN n_22555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.786 122.077 196.814 122.24 ;
      END
   END n_22555

   PIN n_22556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.85 122.077 196.878 122.24 ;
      END
   END n_22556

   PIN n_22569
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 209.65 122.077 209.678 122.24 ;
      END
   END n_22569

   PIN n_22576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.306 122.077 208.334 122.24 ;
      END
   END n_22576

   PIN n_23134
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 222.322 122.077 222.35 122.24 ;
      END
   END n_23134

   PIN n_23144
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.986 122.077 216.014 122.24 ;
      END
   END n_23144

   PIN n_23481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 192.37 122.077 192.398 122.24 ;
      END
   END n_23481

   PIN n_23793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 113.906 241.856 113.934 ;
      END
   END n_23793

   PIN n_23795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 106.098 241.856 106.126 ;
      END
   END n_23795

   PIN n_24123
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 93.746 241.856 93.774 ;
      END
   END n_24123

   PIN n_24149
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 213.874 122.077 213.902 122.24 ;
      END
   END n_24149

   PIN n_24687
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 188.402 122.077 188.43 122.24 ;
      END
   END n_24687

   PIN n_24724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 63.794 241.856 63.822 ;
      END
   END n_24724

   PIN n_24767
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 217.01 122.077 217.038 122.24 ;
      END
   END n_24767

   PIN n_24775
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 118.322 241.856 118.35 ;
      END
   END n_24775

   PIN n_24776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 217.778 122.077 217.806 122.24 ;
      END
   END n_24776

   PIN n_24781
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 63.858 241.856 63.886 ;
      END
   END n_24781

   PIN n_25313
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 213.106 122.077 213.134 122.24 ;
      END
   END n_25313

   PIN n_25456
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 78.322 241.856 78.35 ;
      END
   END n_25456

   PIN n_26039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 219.89 122.077 219.918 122.24 ;
      END
   END n_26039

   PIN n_26051
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 44.594 241.856 44.622 ;
      END
   END n_26051

   PIN n_27859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 77.682 241.856 77.71 ;
      END
   END n_27859

   PIN n_3190
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.258 122.077 110.286 122.24 ;
      END
   END n_3190

   PIN n_32795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.05 122.077 56.078 122.24 ;
      END
   END n_32795

   PIN n_33263
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 29.298 241.856 29.326 ;
      END
   END n_33263

   PIN n_3333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.346 122.077 95.374 122.24 ;
      END
   END n_3333

   PIN n_33852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.794 122.077 127.822 122.24 ;
      END
   END n_33852

   PIN n_34115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.362 122.077 69.39 122.24 ;
      END
   END n_34115

   PIN n_34197
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 171.25 122.077 171.278 122.24 ;
      END
   END n_34197

   PIN n_34198
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.842 122.077 169.87 122.24 ;
      END
   END n_34198

   PIN n_34301
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.41 122.077 39.438 122.24 ;
      END
   END n_34301

   PIN n_34458
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 36.786 241.856 36.814 ;
      END
   END n_34458

   PIN n_34462
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.53 122.077 68.558 122.24 ;
      END
   END n_34462

   PIN n_34463
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.594 122.077 68.622 122.24 ;
      END
   END n_34463

   PIN n_34772
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.042 122.077 53.07 122.24 ;
      END
   END n_34772

   PIN n_34826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 29.17 241.856 29.198 ;
      END
   END n_34826

   PIN n_34941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.586 122.077 65.614 122.24 ;
      END
   END n_34941

   PIN n_35030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 122.077 25.614 122.24 ;
      END
   END n_35030

   PIN n_35071
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 39.858 241.856 39.886 ;
      END
   END n_35071

   PIN n_36024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 29.362 241.856 29.39 ;
      END
   END n_36024

   PIN n_3760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.474 122.077 39.502 122.24 ;
      END
   END n_3760

   PIN n_5402
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.49 122.077 181.518 122.24 ;
      END
   END n_5402

   PIN n_5571
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 166.066 122.077 166.094 122.24 ;
      END
   END n_5571

   PIN n_7597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 75.314 241.856 75.342 ;
      END
   END n_7597

   PIN n_7782
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.954 122.077 115.982 122.24 ;
      END
   END n_7782

   PIN n_7815
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.546 241.856 90.574 ;
      END
   END n_7815

   PIN n_7857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 106.162 241.856 106.19 ;
      END
   END n_7857

   PIN n_9933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 83.314 241.856 83.342 ;
      END
   END n_9933

   PIN FE_OCPN19344_n_142919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 202.034 122.077 202.062 122.24 ;
      END
   END FE_OCPN19344_n_142919

   PIN FE_OFN10229_b_2_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.418 122.077 154.446 122.24 ;
      END
   END FE_OFN10229_b_2_6_2

   PIN FE_OFN10255_b_2_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.514 122.077 150.542 122.24 ;
      END
   END FE_OFN10255_b_2_4_7

   PIN FE_OFN10258_b_2_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.738 122.077 146.766 122.24 ;
      END
   END FE_OFN10258_b_2_4_5

   PIN FE_OFN10270_b_2_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.826 122.077 123.854 122.24 ;
      END
   END FE_OFN10270_b_2_4_1

   PIN FE_OFN10273_b_2_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.098 122.077 162.126 122.24 ;
      END
   END FE_OFN10273_b_2_4_0

   PIN FE_OFN10291_b_2_2_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.698 122.077 123.726 122.24 ;
      END
   END FE_OFN10291_b_2_2_4

   PIN FE_OFN1088_n_20334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 177.65 122.077 177.678 122.24 ;
      END
   END FE_OFN1088_n_20334

   PIN FE_OFN1106_n_19671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 202.098 122.077 202.126 122.24 ;
      END
   END FE_OFN1106_n_19671

   PIN FE_OFN11336_n_143645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.066 122.077 166.094 122.24 ;
      END
   END FE_OFN11336_n_143645

   PIN FE_OFN11351_n_140257
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.89 122.077 115.918 122.24 ;
      END
   END FE_OFN11351_n_140257

   PIN FE_OFN11361_n_143059
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.922 122.077 135.95 122.24 ;
      END
   END FE_OFN11361_n_143059

   PIN FE_OFN11368_n_143045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 168.306 122.077 168.334 122.24 ;
      END
   END FE_OFN11368_n_143045

   PIN FE_OFN11370_n_143045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.906 122.077 113.934 122.24 ;
      END
   END FE_OFN11370_n_143045

   PIN FE_OFN11397_n_140245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.298 122.077 125.326 122.24 ;
      END
   END FE_OFN11397_n_140245

   PIN FE_OFN11427_n_142905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.002 122.077 166.03 122.24 ;
      END
   END FE_OFN11427_n_142905

   PIN FE_OFN11432_n_142919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.018 122.077 204.046 122.24 ;
      END
   END FE_OFN11432_n_142919

   PIN FE_OFN11590_n_143231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.746 122.077 77.774 122.24 ;
      END
   END FE_OFN11590_n_143231

   PIN FE_OFN11596_n_112428
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.778 122.077 81.806 122.24 ;
      END
   END FE_OFN11596_n_112428

   PIN FE_OFN11705_n_142947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 200.562 122.077 200.59 122.24 ;
      END
   END FE_OFN11705_n_142947

   PIN FE_OFN11865_n_143230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.722 122.077 116.75 122.24 ;
      END
   END FE_OFN11865_n_143230

   PIN FE_OFN11869_n_143229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 109.682 241.856 109.71 ;
      END
   END FE_OFN11869_n_143229

   PIN FE_OFN11871_n_143229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.226 122.077 162.254 122.24 ;
      END
   END FE_OFN11871_n_143229

   PIN FE_OFN11875_n_143227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.674 122.077 130.702 122.24 ;
      END
   END FE_OFN11875_n_143227

   PIN FE_OFN11889_n_143104
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.57 122.077 107.598 122.24 ;
      END
   END FE_OFN11889_n_143104

   PIN FE_OFN11896_n_143102
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 154.546 122.077 154.574 122.24 ;
      END
   END FE_OFN11896_n_143102

   PIN FE_OFN11917_n_143048
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.122 122.077 139.15 122.24 ;
      END
   END FE_OFN11917_n_143048

   PIN FE_OFN12298_n_111727
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 102.578 241.856 102.606 ;
      END
   END FE_OFN12298_n_111727

   PIN FE_OFN12309_n_111875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.21 122.158 92.238 122.24 ;
      END
   END FE_OFN12309_n_111875

   PIN FE_OFN12318_n_111878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.722 122.077 100.75 122.24 ;
      END
   END FE_OFN12318_n_111878

   PIN FE_OFN12322_n_112427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.634 122.077 123.662 122.24 ;
      END
   END FE_OFN12322_n_112427

   PIN FE_OFN12325_n_112470
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.162 122.077 98.19 122.24 ;
      END
   END FE_OFN12325_n_112470

   PIN FE_OFN12332_n_137473
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.618 122.077 45.646 122.24 ;
      END
   END FE_OFN12332_n_137473

   PIN FE_OFN12348_n_142991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 83.122 241.856 83.15 ;
      END
   END FE_OFN12348_n_142991

   PIN FE_OFN12350_n_142991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.65 122.077 145.678 122.24 ;
      END
   END FE_OFN12350_n_142991

   PIN FE_OFN12378_n_142908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.994 122.077 123.022 122.24 ;
      END
   END FE_OFN12378_n_142908

   PIN FE_OFN12597_n_111737
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.994 122.077 139.022 122.24 ;
      END
   END FE_OFN12597_n_111737

   PIN FE_OFN12599_n_111738
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.874 122.077 133.902 122.24 ;
      END
   END FE_OFN12599_n_111738

   PIN FE_OFN12609_n_112606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.714 122.158 113.742 122.24 ;
      END
   END FE_OFN12609_n_112606

   PIN FE_OFN12611_n_112608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.666 122.077 127.694 122.24 ;
      END
   END FE_OFN12611_n_112608

   PIN FE_OFN12616_n_112689
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 79.282 241.856 79.31 ;
      END
   END FE_OFN12616_n_112689

   PIN FE_OFN12621_n_112690
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.85 122.077 92.878 122.24 ;
      END
   END FE_OFN12621_n_112690

   PIN FE_OFN12627_n_143646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 135.218 122.077 135.246 122.24 ;
      END
   END FE_OFN12627_n_143646

   PIN FE_OFN12655_n_111913
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.634 241.856 75.662 ;
      END
   END FE_OFN12655_n_111913

   PIN FE_OFN12715_n_142865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 37.106 241.856 37.134 ;
      END
   END FE_OFN12715_n_142865

   PIN FE_OFN12960_n_111998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.774 17.842 241.856 17.87 ;
      END
   END FE_OFN12960_n_111998

   PIN FE_OFN12965_n_112000
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 53.298 241.856 53.326 ;
      END
   END FE_OFN12965_n_112000

   PIN FE_OFN12970_n_112611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 67.506 241.856 67.534 ;
      END
   END FE_OFN12970_n_112611

   PIN FE_OFN12985_n_112681
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 55.858 241.856 55.886 ;
      END
   END FE_OFN12985_n_112681

   PIN FE_OFN13013_n_142950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.77 122.077 158.798 122.24 ;
      END
   END FE_OFN13013_n_142950

   PIN FE_OFN13023_n_142949
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 113.778 241.856 113.806 ;
      END
   END FE_OFN13023_n_142949

   PIN FE_OFN13543_n_143609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 37.362 241.856 37.39 ;
      END
   END FE_OFN13543_n_143609

   PIN FE_OFN13547_n_112256
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 40.882 241.856 40.91 ;
      END
   END FE_OFN13547_n_112256

   PIN FE_OFN13556_n_143397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.794 122.077 135.822 122.24 ;
      END
   END FE_OFN13556_n_143397

   PIN FE_OFN13659_n_112318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 36.85 241.856 36.878 ;
      END
   END FE_OFN13659_n_112318

   PIN FE_OFN13700_n_143384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 17.906 241.856 17.934 ;
      END
   END FE_OFN13700_n_143384

   PIN FE_OFN13708_n_143383
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 45.106 241.856 45.134 ;
      END
   END FE_OFN13708_n_143383

   PIN FE_OFN13818_n_112257
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 34.418 241.856 34.446 ;
      END
   END FE_OFN13818_n_112257

   PIN FE_OFN14269_n_140244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.778 122.077 137.806 122.24 ;
      END
   END FE_OFN14269_n_140244

   PIN FE_OFN14270_n_140244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.114 122.077 112.142 122.24 ;
      END
   END FE_OFN14270_n_140244

   PIN FE_OFN15080_n_19611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 61.042 241.856 61.07 ;
      END
   END FE_OFN15080_n_19611

   PIN FE_OFN15155_n_23384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 98.354 241.856 98.382 ;
      END
   END FE_OFN15155_n_23384

   PIN FE_OFN15251_n_39084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 114.034 241.856 114.062 ;
      END
   END FE_OFN15251_n_39084

   PIN FE_OFN16362_b_2_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 139.314 122.077 139.342 122.24 ;
      END
   END FE_OFN16362_b_2_6_1

   PIN FE_OFN16770_n_16098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 98.482 241.856 98.51 ;
      END
   END FE_OFN16770_n_16098

   PIN FE_OFN16941_n_135332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 36.85 241.856 36.878 ;
      END
   END FE_OFN16941_n_135332

   PIN FE_OFN17141_n_22815
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 94.514 241.856 94.542 ;
      END
   END FE_OFN17141_n_22815

   PIN FE_OFN17145_n_22232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.018 122.077 212.046 122.24 ;
      END
   END FE_OFN17145_n_22232

   PIN FE_OFN17169_n_16270
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 132.85 122.077 132.878 122.24 ;
      END
   END FE_OFN17169_n_16270

   PIN FE_OFN17207_n_21410
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.274 122.077 204.302 122.24 ;
      END
   END FE_OFN17207_n_21410

   PIN FE_OFN17264_n_140245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 118.13 241.856 118.158 ;
      END
   END FE_OFN17264_n_140245

   PIN FE_OFN18602_b_2_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.874 122.077 149.902 122.24 ;
      END
   END FE_OFN18602_b_2_6_0

   PIN FE_OFN18750_n_112550
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.882 122.077 120.91 122.24 ;
      END
   END FE_OFN18750_n_112550

   PIN FE_OFN18809_n_143645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.802 241.856 90.83 ;
      END
   END FE_OFN18809_n_143645

   PIN FE_OFN19061_n_21194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 94.386 241.856 94.414 ;
      END
   END FE_OFN19061_n_21194

   PIN FE_OFN2152_n_19668
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 85.426 241.856 85.454 ;
      END
   END FE_OFN2152_n_19668

   PIN FE_OFN2159_n_19626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 94.514 241.856 94.542 ;
      END
   END FE_OFN2159_n_19626

   PIN FE_OFN2284_n_19629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.826 122.077 155.854 122.24 ;
      END
   END FE_OFN2284_n_19629

   PIN FE_OFN3204_n_14458
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.21 122.077 180.238 122.24 ;
      END
   END FE_OFN3204_n_14458

   PIN FE_OFN3244_n_19948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.762 122.077 155.79 122.24 ;
      END
   END FE_OFN3244_n_19948

   PIN FE_OFN3293_n_8246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 67.634 241.856 67.662 ;
      END
   END FE_OFN3293_n_8246

   PIN FE_OFN3382_n_14610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 44.466 241.856 44.494 ;
      END
   END FE_OFN3382_n_14610

   PIN FE_OFN3441_n_12341
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 118.066 241.856 118.094 ;
      END
   END FE_OFN3441_n_12341

   PIN FE_OFN3505_n_12951
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 135.346 122.077 135.374 122.24 ;
      END
   END FE_OFN3505_n_12951

   PIN FE_OFN3587_n_142906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.194 122.077 110.222 122.24 ;
      END
   END FE_OFN3587_n_142906

   PIN FE_OFN3683_n_142948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.842 122.077 105.87 122.24 ;
      END
   END FE_OFN3683_n_142948

   PIN FE_OFN3701_n_143060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.818 122.077 96.846 122.24 ;
      END
   END FE_OFN3701_n_143060

   PIN FE_OFN3720_n_143241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.058 122.077 139.086 122.24 ;
      END
   END FE_OFN3720_n_143241

   PIN FE_OFN3726_n_143241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.986 122.077 112.014 122.24 ;
      END
   END FE_OFN3726_n_143241

   PIN FE_OFN3737_n_143396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 149.81 122.077 149.838 122.24 ;
      END
   END FE_OFN3737_n_143396

   PIN FE_OFN3743_n_143551
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.57 122.077 123.598 122.24 ;
      END
   END FE_OFN3743_n_143551

   PIN FE_OFN3751_n_143549
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.354 122.077 162.382 122.24 ;
      END
   END FE_OFN3751_n_143549

   PIN FE_OFN596_n_8407
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 101.938 241.856 101.966 ;
      END
   END FE_OFN596_n_8407

   PIN FE_OFN700_n_22202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 88.242 241.856 88.27 ;
      END
   END FE_OFN700_n_22202

   PIN FE_OFN791_n_19612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 240.754 122.077 240.782 122.24 ;
      END
   END FE_OFN791_n_19612

   PIN FE_OFN794_n_20260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.37 122.077 208.398 122.24 ;
      END
   END FE_OFN794_n_20260

   PIN FE_OFN832_n_22177
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 98.418 241.856 98.446 ;
      END
   END FE_OFN832_n_22177

   PIN FE_OFN9231_delay_add_ln34_unr2_unr3_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 71.602 241.856 71.63 ;
      END
   END FE_OFN9231_delay_add_ln34_unr2_unr3_stage2_stallmux_q_15_

   PIN add_5900_51_n_88
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 71.41 241.856 71.438 ;
      END
   END add_5900_51_n_88

   PIN b_0_2_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 37.938 241.856 37.966 ;
      END
   END b_0_2_0

   PIN b_0_2_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 53.618 241.856 53.646 ;
      END
   END b_0_2_1

   PIN b_0_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 32.946 241.856 32.974 ;
      END
   END b_0_2_2

   PIN b_0_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 20.978 241.856 21.006 ;
      END
   END b_0_2_3

   PIN b_0_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 204.786 0.0 204.814 0.082 ;
      END
   END b_0_4_1

   PIN b_0_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 41.138 241.856 41.166 ;
      END
   END b_0_6_0

   PIN b_0_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 44.978 241.856 45.006 ;
      END
   END b_0_6_1

   PIN b_0_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 13.362 241.856 13.39 ;
      END
   END b_0_6_2

   PIN b_0_6_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 234.162 0.0 234.19 0.163 ;
      END
   END b_0_6_5

   PIN b_1_9_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.774 102.706 241.856 102.734 ;
      END
   END b_1_9_0

   PIN b_2_2_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.786 122.077 84.814 122.24 ;
      END
   END b_2_2_0

   PIN b_2_2_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.474 122.077 95.502 122.24 ;
      END
   END b_2_2_1

   PIN b_2_2_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.066 122.077 38.094 122.24 ;
      END
   END b_2_2_11

   PIN b_2_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.698 122.077 107.726 122.24 ;
      END
   END b_2_2_2

   PIN b_2_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.466 122.077 132.494 122.24 ;
      END
   END b_2_2_3

   PIN b_2_2_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.002 122.077 102.03 122.24 ;
      END
   END b_2_2_4

   PIN b_2_2_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.506 122.077 91.534 122.24 ;
      END
   END b_2_2_5

   PIN b_2_2_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.986 122.077 72.014 122.24 ;
      END
   END b_2_2_6

   PIN b_2_2_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.21 122.077 92.238 122.24 ;
      END
   END b_2_2_7

   PIN b_2_2_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.682 122.077 45.71 122.24 ;
      END
   END b_2_2_8

   PIN b_2_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 137.842 122.077 137.87 122.24 ;
      END
   END b_2_4_0

   PIN b_2_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.114 122.077 112.142 122.24 ;
      END
   END b_2_4_1

   PIN b_2_4_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.938 122.077 133.966 122.24 ;
      END
   END b_2_4_11

   PIN b_2_4_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.562 122.077 112.59 122.24 ;
      END
   END b_2_4_12

   PIN b_2_4_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.234 122.077 101.262 122.24 ;
      END
   END b_2_4_13

   PIN b_2_4_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.362 122.077 101.39 122.24 ;
      END
   END b_2_4_2

   PIN b_2_4_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 137.138 122.077 137.166 122.24 ;
      END
   END b_2_4_3

   PIN b_2_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 132.914 122.077 132.942 122.24 ;
      END
   END b_2_4_4

   PIN b_2_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.346 122.077 79.374 122.24 ;
      END
   END b_2_4_5

   PIN b_2_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.058 122.077 91.086 122.24 ;
      END
   END b_2_4_6

   PIN b_2_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.786 122.077 116.814 122.24 ;
      END
   END b_2_4_7

   PIN b_2_4_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.738 122.077 106.766 122.24 ;
      END
   END b_2_4_8

   PIN b_2_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 129.01 122.077 129.038 122.24 ;
      END
   END b_2_6_1

   PIN b_2_6_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.738 122.077 130.766 122.24 ;
      END
   END b_2_6_10

   PIN b_2_6_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.97 122.077 113.998 122.24 ;
      END
   END b_2_6_11

   PIN b_2_6_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.93 122.077 122.958 122.24 ;
      END
   END b_2_6_12

   PIN b_2_6_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.842 122.077 113.87 122.24 ;
      END
   END b_2_6_13

   PIN b_2_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 125.042 122.077 125.07 122.24 ;
      END
   END b_2_6_2

   PIN b_2_6_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.714 122.077 145.742 122.24 ;
      END
   END b_2_6_3

   PIN b_2_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.674 122.077 146.702 122.24 ;
      END
   END b_2_6_4

   PIN b_2_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.642 122.077 150.67 122.24 ;
      END
   END b_2_6_7

   PIN b_2_6_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 118.386 122.077 118.414 122.24 ;
      END
   END b_2_6_9

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 212.146 122.158 212.174 122.24 ;
      END
   END ispd_clk

   PIN mul_4370_72_n_149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 37.042 241.856 37.07 ;
      END
   END mul_4370_72_n_149

   PIN mul_4370_72_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 4.85 241.856 4.878 ;
      END
   END mul_4370_72_n_50

   PIN mul_4370_72_n_66
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 4.786 241.856 4.814 ;
      END
   END mul_4370_72_n_66

   PIN mul_4370_72_n_793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 2.354 241.856 2.382 ;
      END
   END mul_4370_72_n_793

   PIN mul_4370_72_n_840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 20.786 241.856 20.814 ;
      END
   END mul_4370_72_n_840

   PIN mul_4377_72_n_106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 83.378 241.856 83.406 ;
      END
   END mul_4377_72_n_106

   PIN mul_4377_72_n_114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 71.666 241.856 71.694 ;
      END
   END mul_4377_72_n_114

   PIN mul_4377_72_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.994 241.856 91.022 ;
      END
   END mul_4377_72_n_116

   PIN mul_4665_72_n_244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.794 122.077 119.822 122.24 ;
      END
   END mul_4665_72_n_244

   PIN mul_4665_72_n_330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.226 122.077 66.254 122.24 ;
      END
   END mul_4665_72_n_330

   PIN mul_4665_72_n_338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.106 122.077 13.134 122.24 ;
      END
   END mul_4665_72_n_338

   PIN mul_4665_72_n_339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.962 122.077 6.99 122.24 ;
      END
   END mul_4665_72_n_339

   PIN mul_4667_72_n_334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.338 122.077 100.366 122.24 ;
      END
   END mul_4667_72_n_334

   PIN mul_4667_72_n_340
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.946 122.077 96.974 122.24 ;
      END
   END mul_4667_72_n_340

   PIN mul_4669_72_n_315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.81 122.077 117.838 122.24 ;
      END
   END mul_4669_72_n_315

   PIN mul_4669_72_n_340
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 140.85 122.077 140.878 122.24 ;
      END
   END mul_4669_72_n_340

   PIN mul_ln34_unr2_unr2_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.29 122.077 66.318 122.24 ;
      END
   END mul_ln34_unr2_unr2_z_11_

   PIN mul_ln34_unr2_unr5_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 40.818 241.856 40.846 ;
      END
   END mul_ln34_unr2_unr5_z_13_

   PIN mul_ln34_unr2_unr5_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 45.17 241.856 45.198 ;
      END
   END mul_ln34_unr2_unr5_z_14_

   PIN n_10106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.33 122.077 89.358 122.24 ;
      END
   END n_10106

   PIN n_10396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.034 122.077 106.062 122.24 ;
      END
   END n_10396

   PIN n_10648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 113.97 241.856 113.998 ;
      END
   END n_10648

   PIN n_10996
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 13.618 241.856 13.646 ;
      END
   END n_10996

   PIN n_10998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 55.794 241.856 55.822 ;
      END
   END n_10998

   PIN n_111930
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 53.298 241.856 53.326 ;
      END
   END n_111930

   PIN n_112180
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.018 122.077 76.046 122.24 ;
      END
   END n_112180

   PIN n_112566
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.642 122.077 86.67 122.24 ;
      END
   END n_112566

   PIN n_112607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.21 122.158 116.238 122.24 ;
      END
   END n_112607

   PIN n_112707
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.738 241.856 90.766 ;
      END
   END n_112707

   PIN n_112826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.098 122.077 66.126 122.24 ;
      END
   END n_112826

   PIN n_112827
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.034 122.077 66.062 122.24 ;
      END
   END n_112827

   PIN n_112875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.354 122.077 66.382 122.24 ;
      END
   END n_112875

   PIN n_112887
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 44.402 241.856 44.43 ;
      END
   END n_112887

   PIN n_112910
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.458 241.856 25.486 ;
      END
   END n_112910

   PIN n_112911
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.586 241.856 25.614 ;
      END
   END n_112911

   PIN n_112930
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 29.042 241.856 29.07 ;
      END
   END n_112930

   PIN n_113050
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 32.178 241.856 32.206 ;
      END
   END n_113050

   PIN n_113218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.946 122.077 96.974 122.24 ;
      END
   END n_113218

   PIN n_113364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 52.018 241.856 52.046 ;
      END
   END n_113364

   PIN n_113365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 54.578 241.856 54.606 ;
      END
   END n_113365

   PIN n_113366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 40.562 241.856 40.59 ;
      END
   END n_113366

   PIN n_113426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 48.498 241.856 48.526 ;
      END
   END n_113426

   PIN n_113502
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.658 122.077 92.686 122.24 ;
      END
   END n_113502

   PIN n_113544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.906 122.077 169.934 122.24 ;
      END
   END n_113544

   PIN n_113546
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.154 122.077 135.182 122.24 ;
      END
   END n_113546

   PIN n_113561
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.258 122.077 158.286 122.24 ;
      END
   END n_113561

   PIN n_113602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 44.338 241.856 44.366 ;
      END
   END n_113602

   PIN n_113603
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 45.234 241.856 45.262 ;
      END
   END n_113603

   PIN n_113699
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.274 122.077 140.302 122.24 ;
      END
   END n_113699

   PIN n_113855
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.722 122.077 92.75 122.24 ;
      END
   END n_113855

   PIN n_113856
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.45 122.077 94.478 122.24 ;
      END
   END n_113856

   PIN n_113866
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.89 122.077 67.918 122.24 ;
      END
   END n_113866

   PIN n_113926
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.202 122.077 113.23 122.24 ;
      END
   END n_113926

   PIN n_113994
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.674 122.077 18.702 122.24 ;
      END
   END n_113994

   PIN n_114084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.978 122.077 37.006 122.24 ;
      END
   END n_114084

   PIN n_114198
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.97 122.077 65.998 122.24 ;
      END
   END n_114198

   PIN n_114263
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.754 122.077 96.782 122.24 ;
      END
   END n_114263

   PIN n_114274
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.754 122.077 56.782 122.24 ;
      END
   END n_114274

   PIN n_114292
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 34.482 241.856 34.51 ;
      END
   END n_114292

   PIN n_114416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.338 122.077 140.366 122.24 ;
      END
   END n_114416

   PIN n_114432
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.922 122.077 119.95 122.24 ;
      END
   END n_114432

   PIN n_114581
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 21.17 241.856 21.198 ;
      END
   END n_114581

   PIN n_114701
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.77 122.077 94.798 122.24 ;
      END
   END n_114701

   PIN n_115305
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.762 122.077 147.79 122.24 ;
      END
   END n_115305

   PIN n_11535
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.906 122.077 105.934 122.24 ;
      END
   END n_11535

   PIN n_115461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.042 122.077 37.07 122.24 ;
      END
   END n_115461

   PIN n_115480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.042 122.077 109.07 122.24 ;
      END
   END n_115480

   PIN n_115635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.178 122.077 112.206 122.24 ;
      END
   END n_115635

   PIN n_115636
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.05 122.077 112.078 122.24 ;
      END
   END n_115636

   PIN n_116469
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.37 122.077 112.398 122.24 ;
      END
   END n_116469

   PIN n_117228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 71.538 241.856 71.566 ;
      END
   END n_117228

   PIN n_117236
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 94.578 241.856 94.606 ;
      END
   END n_117236

   PIN n_117237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 94.258 241.856 94.286 ;
      END
   END n_117237

   PIN n_117368
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.362 122.077 117.39 122.24 ;
      END
   END n_117368

   PIN n_117402
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 71.346 241.856 71.374 ;
      END
   END n_117402

   PIN n_117521
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.226 122.077 66.254 122.24 ;
      END
   END n_117521

   PIN n_118323
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.386 122.077 62.414 122.24 ;
      END
   END n_118323

   PIN n_119297
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.082 122.077 84.11 122.24 ;
      END
   END n_119297

   PIN n_119298
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.826 122.077 83.854 122.24 ;
      END
   END n_119298

   PIN n_119316
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.746 122.077 109.774 122.24 ;
      END
   END n_119316

   PIN n_119738
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.258 122.077 62.286 122.24 ;
      END
   END n_119738

   PIN n_119899
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 79.538 241.856 79.566 ;
      END
   END n_119899

   PIN n_119933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 53.426 241.856 53.454 ;
      END
   END n_119933

   PIN n_119934
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 53.362 241.856 53.39 ;
      END
   END n_119934

   PIN n_119959
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 40.754 241.856 40.782 ;
      END
   END n_119959

   PIN n_119983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.746 122.077 45.774 122.24 ;
      END
   END n_119983

   PIN n_120078
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.642 122.077 94.67 122.24 ;
      END
   END n_120078

   PIN n_120079
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.298 122.077 93.326 122.24 ;
      END
   END n_120079

   PIN n_120193
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 56.37 241.856 56.398 ;
      END
   END n_120193

   PIN n_120437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 75.378 241.856 75.406 ;
      END
   END n_120437

   PIN n_120635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.322 122.077 94.35 122.24 ;
      END
   END n_120635

   PIN n_120746
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.962 122.077 134.99 122.24 ;
      END
   END n_120746

   PIN n_120996
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.602 122.077 55.63 122.24 ;
      END
   END n_120996

   PIN n_121285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 78.898 241.856 78.926 ;
      END
   END n_121285

   PIN n_121633
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 87.218 241.856 87.246 ;
      END
   END n_121633

   PIN n_121772
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.522 122.077 81.55 122.24 ;
      END
   END n_121772

   PIN n_121803
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 17.65 241.856 17.678 ;
      END
   END n_121803

   PIN n_121832
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 13.106 241.856 13.134 ;
      END
   END n_121832

   PIN n_121834
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 13.234 241.856 13.262 ;
      END
   END n_121834

   PIN n_121906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.93 122.077 138.958 122.24 ;
      END
   END n_121906

   PIN n_121932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 86.578 241.856 86.606 ;
      END
   END n_121932

   PIN n_121933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 86.642 241.856 86.67 ;
      END
   END n_121933

   PIN n_122107
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.746 122.077 5.774 122.24 ;
      END
   END n_122107

   PIN n_122555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 36.978 241.856 37.006 ;
      END
   END n_122555

   PIN n_122556
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 48.178 241.856 48.206 ;
      END
   END n_122556

   PIN n_12342
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 117.618 241.856 117.646 ;
      END
   END n_12342

   PIN n_123546
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 4.658 241.856 4.686 ;
      END
   END n_123546

   PIN n_123558
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 17.586 241.856 17.614 ;
      END
   END n_123558

   PIN n_123606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.93 122.077 50.958 122.24 ;
      END
   END n_123606

   PIN n_123620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 20.722 241.856 20.75 ;
      END
   END n_123620

   PIN n_123678
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.162 122.077 162.19 122.24 ;
      END
   END n_123678

   PIN n_123759
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.394 241.856 25.422 ;
      END
   END n_123759

   PIN n_124048
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.962 122.077 142.99 122.24 ;
      END
   END n_124048

   PIN n_124617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.898 122.077 142.926 122.24 ;
      END
   END n_124617

   PIN n_124974
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.802 122.077 130.83 122.24 ;
      END
   END n_124974

   PIN n_124975
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.866 122.077 130.894 122.24 ;
      END
   END n_124975

   PIN n_125043
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 69.49 241.856 69.518 ;
      END
   END n_125043

   PIN n_125044
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 67.378 241.856 67.406 ;
      END
   END n_125044

   PIN n_125081
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 93.682 241.856 93.71 ;
      END
   END n_125081

   PIN n_125082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 88.178 241.856 88.206 ;
      END
   END n_125082

   PIN n_125769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 13.042 241.856 13.07 ;
      END
   END n_125769

   PIN n_125781
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 13.042 241.856 13.07 ;
      END
   END n_125781

   PIN n_125786
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 12.978 241.856 13.006 ;
      END
   END n_125786

   PIN n_12587
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.018 122.077 116.046 122.24 ;
      END
   END n_12587

   PIN n_126291
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 59.89 241.856 59.918 ;
      END
   END n_126291

   PIN n_126292
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 69.426 241.856 69.454 ;
      END
   END n_126292

   PIN n_126559
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 17.842 241.856 17.87 ;
      END
   END n_126559

   PIN n_126560
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 17.778 241.856 17.806 ;
      END
   END n_126560

   PIN n_12711
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.25 241.856 75.278 ;
      END
   END n_12711

   PIN n_127736
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 71.218 241.856 71.246 ;
      END
   END n_127736

   PIN n_127873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 9.906 241.856 9.934 ;
      END
   END n_127873

   PIN n_127889
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.69 122.077 48.718 122.24 ;
      END
   END n_127889

   PIN n_127896
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 33.074 241.856 33.102 ;
      END
   END n_127896

   PIN n_127954
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 21.298 241.856 21.326 ;
      END
   END n_127954

   PIN n_128003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.826 122.077 27.854 122.24 ;
      END
   END n_128003

   PIN n_128515
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 59.826 241.856 59.854 ;
      END
   END n_128515

   PIN n_128527
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 61.618 241.856 61.646 ;
      END
   END n_128527

   PIN n_128971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.594 122.077 36.622 122.24 ;
      END
   END n_128971

   PIN n_128973
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.53 122.077 36.558 122.24 ;
      END
   END n_128973

   PIN n_129101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.538 122.077 127.566 122.24 ;
      END
   END n_129101

   PIN n_12956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.818 122.077 120.846 122.24 ;
      END
   END n_12956

   PIN n_130212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.29 122.077 34.318 122.24 ;
      END
   END n_130212

   PIN n_130734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.954 122.077 123.982 122.24 ;
      END
   END n_130734

   PIN n_131017
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.346 122.077 39.374 122.24 ;
      END
   END n_131017

   PIN n_131069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 72.69 122.077 72.718 122.24 ;
      END
   END n_131069

   PIN n_131070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.562 122.077 72.59 122.24 ;
      END
   END n_131070

   PIN n_131430
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.29 122.077 66.318 122.24 ;
      END
   END n_131430

   PIN n_131641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.714 122.077 81.742 122.24 ;
      END
   END n_131641

   PIN n_132252
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.218 122.077 103.246 122.24 ;
      END
   END n_132252

   PIN n_132417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 29.234 241.856 29.262 ;
      END
   END n_132417

   PIN n_132434
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 36.722 241.856 36.75 ;
      END
   END n_132434

   PIN n_132699
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.538 122.077 55.566 122.24 ;
      END
   END n_132699

   PIN n_132892
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.586 122.077 57.614 122.24 ;
      END
   END n_132892

   PIN n_132893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.522 122.077 57.55 122.24 ;
      END
   END n_132893

   PIN n_132961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.714 122.077 73.742 122.24 ;
      END
   END n_132961

   PIN n_132962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.522 122.077 73.55 122.24 ;
      END
   END n_132962

   PIN n_133201
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.194 122.077 62.222 122.24 ;
      END
   END n_133201

   PIN n_133273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 136.05 122.077 136.078 122.24 ;
      END
   END n_133273

   PIN n_133287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.77 122.077 142.798 122.24 ;
      END
   END n_133287

   PIN n_133303
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.794 122.077 103.822 122.24 ;
      END
   END n_133303

   PIN n_133427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.834 122.077 142.862 122.24 ;
      END
   END n_133427

   PIN n_133450
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 29.106 241.856 29.134 ;
      END
   END n_133450

   PIN n_133506
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.338 122.077 132.366 122.24 ;
      END
   END n_133506

   PIN n_133858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 36.658 241.856 36.686 ;
      END
   END n_133858

   PIN n_133861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.81 122.077 69.838 122.24 ;
      END
   END n_133861

   PIN n_133939
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.202 241.856 25.23 ;
      END
   END n_133939

   PIN n_134000
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.938 122.077 69.966 122.24 ;
      END
   END n_134000

   PIN n_134256
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.138 241.856 25.166 ;
      END
   END n_134256

   PIN n_134400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.434 122.077 104.462 122.24 ;
      END
   END n_134400

   PIN n_134706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 30.002 241.856 30.03 ;
      END
   END n_134706

   PIN n_134708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 56.818 241.856 56.846 ;
      END
   END n_134708

   PIN n_134825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 135.858 122.077 135.886 122.24 ;
      END
   END n_134825

   PIN n_134924
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.874 122.077 69.902 122.24 ;
      END
   END n_134924

   PIN n_134992
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.026 122.077 47.054 122.24 ;
      END
   END n_134992

   PIN n_135296
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 21.362 241.856 21.39 ;
      END
   END n_135296

   PIN n_135308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.858 122.077 135.886 122.24 ;
      END
   END n_135308

   PIN n_135370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 82.674 241.856 82.702 ;
      END
   END n_135370

   PIN n_135438
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.762 122.077 123.79 122.24 ;
      END
   END n_135438

   PIN n_135524
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.282 122.077 39.31 122.24 ;
      END
   END n_135524

   PIN n_135528
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.338 122.077 108.366 122.24 ;
      END
   END n_135528

   PIN n_135704
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 20.85 241.856 20.878 ;
      END
   END n_135704

   PIN n_135859
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.882 122.077 8.91 122.24 ;
      END
   END n_135859

   PIN n_135947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.546 122.077 58.574 122.24 ;
      END
   END n_135947

   PIN n_135957
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.05 122.077 56.078 122.24 ;
      END
   END n_135957

   PIN n_136054
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 28.978 241.856 29.006 ;
      END
   END n_136054

   PIN n_136077
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 12.466 241.856 12.494 ;
      END
   END n_136077

   PIN n_136078
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 10.226 241.856 10.254 ;
      END
   END n_136078

   PIN n_136095
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 165.362 122.077 165.39 122.24 ;
      END
   END n_136095

   PIN n_136295
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 21.298 241.856 21.326 ;
      END
   END n_136295

   PIN n_136526
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.81 122.077 53.838 122.24 ;
      END
   END n_136526

   PIN n_136551
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 12.402 241.856 12.43 ;
      END
   END n_136551

   PIN n_136552
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 10.162 241.856 10.19 ;
      END
   END n_136552

   PIN n_136555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 12.338 241.856 12.366 ;
      END
   END n_136555

   PIN n_136727
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 4.658 241.856 4.686 ;
      END
   END n_136727

   PIN n_136754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 10.098 241.856 10.126 ;
      END
   END n_136754

   PIN n_136800
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 25.266 241.856 25.294 ;
      END
   END n_136800

   PIN n_136807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.186 241.856 75.214 ;
      END
   END n_136807

   PIN n_136808
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 85.298 241.856 85.326 ;
      END
   END n_136808

   PIN n_136922
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 177.458 122.077 177.486 122.24 ;
      END
   END n_136922

   PIN n_136951
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 63.602 241.856 63.63 ;
      END
   END n_136951

   PIN n_137637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.746 122.077 53.774 122.24 ;
      END
   END n_137637

   PIN n_137650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 10.034 241.856 10.062 ;
      END
   END n_137650

   PIN n_14254
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.122 122.077 131.15 122.24 ;
      END
   END n_14254

   PIN n_14255
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 131.442 122.077 131.47 122.24 ;
      END
   END n_14255

   PIN n_14287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 127.666 122.077 127.694 122.24 ;
      END
   END n_14287

   PIN n_142906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 109.746 241.856 109.774 ;
      END
   END n_142906

   PIN n_142909
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 110.002 241.856 110.03 ;
      END
   END n_142909

   PIN n_143255
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 13.17 241.856 13.198 ;
      END
   END n_143255

   PIN n_143341
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 40.818 241.856 40.846 ;
      END
   END n_143341

   PIN n_143721
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.874 122.077 77.902 122.24 ;
      END
   END n_143721

   PIN n_143848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.25 122.077 43.278 122.24 ;
      END
   END n_143848

   PIN n_144235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 102.002 241.856 102.03 ;
      END
   END n_144235

   PIN n_144239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 117.554 241.856 117.582 ;
      END
   END n_144239

   PIN n_144318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 60.018 241.856 60.046 ;
      END
   END n_144318

   PIN n_14452
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 63.666 241.856 63.694 ;
      END
   END n_14452

   PIN n_14557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 98.29 241.856 98.318 ;
      END
   END n_14557

   PIN n_14659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.506 122.077 227.534 122.24 ;
      END
   END n_14659

   PIN n_14956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.082 122.077 212.11 122.24 ;
      END
   END n_14956

   PIN n_15206
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 98.226 241.856 98.254 ;
      END
   END n_15206

   PIN n_15462
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.954 122.077 211.982 122.24 ;
      END
   END n_15462

   PIN n_16034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 102.066 241.856 102.094 ;
      END
   END n_16034

   PIN n_16166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 177.586 122.077 177.614 122.24 ;
      END
   END n_16166

   PIN n_16255
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 40.69 241.856 40.718 ;
      END
   END n_16255

   PIN n_16364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 86.706 241.856 86.734 ;
      END
   END n_16364

   PIN n_16366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 9.97 241.856 9.998 ;
      END
   END n_16366

   PIN n_16486
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 105.906 241.856 105.934 ;
      END
   END n_16486

   PIN n_17494
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.418 241.856 90.446 ;
      END
   END n_17494

   PIN n_17661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 118.45 241.856 118.478 ;
      END
   END n_17661

   PIN n_17796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 106.098 241.856 106.126 ;
      END
   END n_17796

   PIN n_18022
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 110.322 241.856 110.35 ;
      END
   END n_18022

   PIN n_18128
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 12.978 241.856 13.006 ;
      END
   END n_18128

   PIN n_18199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.442 122.077 227.47 122.24 ;
      END
   END n_18199

   PIN n_18869
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 67.634 241.856 67.662 ;
      END
   END n_18869

   PIN n_18877
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 59.954 241.856 59.982 ;
      END
   END n_18877

   PIN n_18948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 20.658 241.856 20.686 ;
      END
   END n_18948

   PIN n_18989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 101.938 241.856 101.966 ;
      END
   END n_18989

   PIN n_19350
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.282 122.077 231.31 122.24 ;
      END
   END n_19350

   PIN n_19373
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.858 122.077 215.886 122.24 ;
      END
   END n_19373

   PIN n_19607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 48.562 241.856 48.59 ;
      END
   END n_19607

   PIN n_19629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 86.77 241.856 86.798 ;
      END
   END n_19629

   PIN n_19657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 63.794 241.856 63.822 ;
      END
   END n_19657

   PIN n_19681
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 83.058 241.856 83.086 ;
      END
   END n_19681

   PIN n_19914
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 44.53 241.856 44.558 ;
      END
   END n_19914

   PIN n_19971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 63.922 241.856 63.95 ;
      END
   END n_19971

   PIN n_19983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 98.61 241.856 98.638 ;
      END
   END n_19983

   PIN n_20006
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 60.082 241.856 60.11 ;
      END
   END n_20006

   PIN n_20085
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 82.994 241.856 83.022 ;
      END
   END n_20085

   PIN n_20090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 82.93 241.856 82.958 ;
      END
   END n_20090

   PIN n_20275
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 17.714 241.856 17.742 ;
      END
   END n_20275

   PIN n_20413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.634 122.077 155.662 122.24 ;
      END
   END n_20413

   PIN n_20639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 79.218 241.856 79.246 ;
      END
   END n_20639

   PIN n_20872
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 56.306 241.856 56.334 ;
      END
   END n_20872

   PIN n_21109
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 79.154 241.856 79.182 ;
      END
   END n_21109

   PIN n_21129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 98.354 241.856 98.382 ;
      END
   END n_21129

   PIN n_21187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 110.258 241.856 110.286 ;
      END
   END n_21187

   PIN n_21414
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 94.642 241.856 94.67 ;
      END
   END n_21414

   PIN n_21637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 56.178 241.856 56.206 ;
      END
   END n_21637

   PIN n_21657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 59.762 241.856 59.79 ;
      END
   END n_21657

   PIN n_21680
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 94.45 241.856 94.478 ;
      END
   END n_21680

   PIN n_21703
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 118.002 241.856 118.03 ;
      END
   END n_21703

   PIN n_21708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 75.57 241.856 75.598 ;
      END
   END n_21708

   PIN n_21709
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.93 241.856 90.958 ;
      END
   END n_21709

   PIN n_21771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.73 122.077 71.758 122.24 ;
      END
   END n_21771

   PIN n_21806
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.858 122.077 71.886 122.24 ;
      END
   END n_21806

   PIN n_22159
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.922 122.077 71.95 122.24 ;
      END
   END n_22159

   PIN n_22224
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 118.386 241.856 118.414 ;
      END
   END n_22224

   PIN n_22231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.674 241.856 90.702 ;
      END
   END n_22231

   PIN n_22243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 79.09 241.856 79.118 ;
      END
   END n_22243

   PIN n_22795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 113.714 241.856 113.742 ;
      END
   END n_22795

   PIN n_22822
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 79.026 241.856 79.054 ;
      END
   END n_22822

   PIN n_23394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 90.738 241.856 90.766 ;
      END
   END n_23394

   PIN n_23404
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 79.218 241.856 79.246 ;
      END
   END n_23404

   PIN n_23460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 193.01 122.077 193.038 122.24 ;
      END
   END n_23460

   PIN n_24014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 52.21 241.856 52.238 ;
      END
   END n_24014

   PIN n_24074
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 109.618 241.856 109.646 ;
      END
   END n_24074

   PIN n_24124
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 217.266 122.077 217.294 122.24 ;
      END
   END n_24124

   PIN n_24141
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 93.618 241.856 93.646 ;
      END
   END n_24141

   PIN n_24645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 40.69 241.856 40.718 ;
      END
   END n_24645

   PIN n_24723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 48.498 241.856 48.526 ;
      END
   END n_24723

   PIN n_24774
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 117.938 241.856 117.966 ;
      END
   END n_24774

   PIN n_25460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 85.618 241.856 85.646 ;
      END
   END n_25460

   PIN n_26642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 83.698 241.856 83.726 ;
      END
   END n_26642

   PIN n_28886
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 90.61 241.856 90.638 ;
      END
   END n_28886

   PIN n_31620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.178 122.077 96.206 122.24 ;
      END
   END n_31620

   PIN n_31789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 36.914 241.856 36.942 ;
      END
   END n_31789

   PIN n_32482
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 33.266 241.856 33.294 ;
      END
   END n_32482

   PIN n_32483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 33.202 241.856 33.23 ;
      END
   END n_32483

   PIN n_32637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.314 122.077 131.342 122.24 ;
      END
   END n_32637

   PIN n_32919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.242 122.077 16.27 122.24 ;
      END
   END n_32919

   PIN n_32920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.498 122.077 16.526 122.24 ;
      END
   END n_32920

   PIN n_32934
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.762 122.077 27.79 122.24 ;
      END
   END n_32934

   PIN n_33003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.25 122.077 43.278 122.24 ;
      END
   END n_33003

   PIN n_33076
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.17 122.077 133.198 122.24 ;
      END
   END n_33076

   PIN n_33077
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.602 122.077 127.63 122.24 ;
      END
   END n_33077

   PIN n_33264
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 25.522 241.856 25.55 ;
      END
   END n_33264

   PIN n_33268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 29.938 241.856 29.966 ;
      END
   END n_33268

   PIN n_33473
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.506 122.077 123.534 122.24 ;
      END
   END n_33473

   PIN n_33483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.746 122.077 69.774 122.24 ;
      END
   END n_33483

   PIN n_33921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.89 122.077 27.918 122.24 ;
      END
   END n_33921

   PIN n_33953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.106 122.077 53.134 122.24 ;
      END
   END n_33953

   PIN n_34366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.858 122.077 47.886 122.24 ;
      END
   END n_34366

   PIN n_34708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 173.682 122.077 173.71 122.24 ;
      END
   END n_34708

   PIN n_34720
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 127.73 122.077 127.758 122.24 ;
      END
   END n_34720

   PIN n_35010
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.274 122.077 108.302 122.24 ;
      END
   END n_35010

   PIN n_35016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.45 122.077 54.478 122.24 ;
      END
   END n_35016

   PIN n_35029
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.778 122.077 25.806 122.24 ;
      END
   END n_35029

   PIN n_35032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.61 122.077 26.638 122.24 ;
      END
   END n_35032

   PIN n_35033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.306 122.077 56.334 122.24 ;
      END
   END n_35033

   PIN n_35070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 29.426 241.856 29.454 ;
      END
   END n_35070

   PIN n_35739
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.746 122.077 117.774 122.24 ;
      END
   END n_35739

   PIN n_36449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.09 122.077 135.118 122.24 ;
      END
   END n_36449

   PIN n_3711
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.21 122.077 84.238 122.24 ;
      END
   END n_3711

   PIN n_3868
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.93 122.077 130.958 122.24 ;
      END
   END n_3868

   PIN n_39087
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.362 122.077 181.39 122.24 ;
      END
   END n_39087

   PIN n_39278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.858 122.077 119.886 122.24 ;
      END
   END n_39278

   PIN n_3945
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 4.722 241.856 4.75 ;
      END
   END n_3945

   PIN n_39484
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.986 122.077 112.014 122.24 ;
      END
   END n_39484

   PIN n_39485
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.05 122.077 112.078 122.24 ;
      END
   END n_39485

   PIN n_41711
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 241.693 68.85 241.856 68.878 ;
      END
   END n_41711

   PIN n_4199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.002 122.077 70.03 122.24 ;
      END
   END n_4199

   PIN n_5193
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.618 122.077 77.646 122.24 ;
      END
   END n_5193

   PIN n_5196
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.018 122.077 84.046 122.24 ;
      END
   END n_5196

   PIN n_5565
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.65 122.077 81.678 122.24 ;
      END
   END n_5565

   PIN n_6522
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.402 122.077 132.43 122.24 ;
      END
   END n_6522

   PIN n_6525
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.762 122.077 123.79 122.24 ;
      END
   END n_6525

   PIN n_6542
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.802 122.077 106.83 122.24 ;
      END
   END n_6542

   PIN n_6619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.098 122.077 106.126 122.24 ;
      END
   END n_6619

   PIN n_6693
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.05 122.077 120.078 122.24 ;
      END
   END n_6693

   PIN n_6697
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.082 122.077 116.11 122.24 ;
      END
   END n_6697

   PIN n_6937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 63.986 241.856 64.014 ;
      END
   END n_6937

   PIN n_7273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 40.498 241.856 40.526 ;
      END
   END n_7273

   PIN n_8119
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.866 122.077 50.894 122.24 ;
      END
   END n_8119

   PIN n_8247
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 62.898 241.856 62.926 ;
      END
   END n_8247

   PIN n_8343
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 52.146 241.856 52.174 ;
      END
   END n_8343

   PIN n_8387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 78.258 241.856 78.286 ;
      END
   END n_8387

   PIN n_890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 150.642 122.077 150.67 122.24 ;
      END
   END n_890

   PIN n_912
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 241.693 109.938 241.856 109.966 ;
      END
   END n_912

   PIN n_9132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.146 122.077 212.174 122.24 ;
      END
   END n_9132

   PIN n_9798
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.85 122.077 140.878 122.24 ;
      END
   END n_9798

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 241.856 122.24 ;
      LAYER V1 ;
         RECT 0.0 0.0 241.856 122.24 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 241.856 122.24 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 241.856 122.24 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 241.856 122.24 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 241.856 122.24 ;
      LAYER M1 ;
         RECT 0.0 0.0 241.856 122.24 ;
   END
END h0_mgc_matrix_mult_a

MACRO h9_mgc_matrix_mult_b
   CLASS BLOCK ;
   FOREIGN h9 ;
   ORIGIN 0 0 ;
   SIZE 85.568 BY 75.53 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1072_n_16034
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.41 0.0 31.438 0.163 ;
      END
   END FE_OFN1072_n_16034

   PIN FE_OFN12071_n_41544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.282 75.366 23.31 75.529 ;
      END
   END FE_OFN12071_n_41544

   PIN FE_OFN12072_n_41544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 71.986 0.163 72.014 ;
      END
   END FE_OFN12072_n_41544

   PIN FE_OFN13275_n_143160
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.114 75.366 24.142 75.529 ;
      END
   END FE_OFN13275_n_143160

   PIN FE_OFN13371_n_41505
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.458 75.366 25.486 75.529 ;
      END
   END FE_OFN13371_n_41505

   PIN FE_OFN13374_n_41505
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.074 75.366 17.102 75.529 ;
      END
   END FE_OFN13374_n_41505

   PIN FE_OFN13923_n_143215
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.114 0.163 72.142 ;
      END
   END FE_OFN13923_n_143215

   PIN FE_OFN13929_n_143214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 61.106 0.163 61.134 ;
      END
   END FE_OFN13929_n_143214

   PIN FE_OFN13930_n_143214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.37 75.366 8.398 75.529 ;
      END
   END FE_OFN13930_n_143214

   PIN FE_OFN13940_n_143187
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.21 0.163 68.238 ;
      END
   END FE_OFN13940_n_143187

   PIN FE_OFN13972_n_41362
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.562 0.163 72.59 ;
      END
   END FE_OFN13972_n_41362

   PIN FE_OFN13973_n_41362
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.01 75.366 17.038 75.529 ;
      END
   END FE_OFN13973_n_41362

   PIN FE_OFN14504_n_41536
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 65.394 0.163 65.422 ;
      END
   END FE_OFN14504_n_41536

   PIN FE_OFN14973_n_67017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.722 0.0 4.75 0.163 ;
      END
   END FE_OFN14973_n_67017

   PIN FE_OFN17078_n_140296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.474 75.366 55.502 75.529 ;
      END
   END FE_OFN17078_n_140296

   PIN FE_OFN17700_delay_mul_ln34_unr6_unr8_stage2_stallmux_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.226 75.366 42.254 75.529 ;
      END
   END FE_OFN17700_delay_mul_ln34_unr6_unr8_stage2_stallmux_z_2_

   PIN FE_OFN18514_delay_add_ln34_unr2_unr2_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.362 0.163 29.39 ;
      END
   END FE_OFN18514_delay_add_ln34_unr2_unr2_stage2_stallmux_q_13_

   PIN FE_OFN5666_delay_mul_ln34_unr6_unr3_stage2_stallmux_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 48.562 85.568 48.59 ;
      END
   END FE_OFN5666_delay_mul_ln34_unr6_unr3_stage2_stallmux_z_2_

   PIN FE_OFN5813_delay_mul_ln34_unr6_unr4_stage2_stallmux_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 60.146 85.568 60.174 ;
      END
   END FE_OFN5813_delay_mul_ln34_unr6_unr4_stage2_stallmux_z_2_

   PIN FE_OFN5889_n_41535
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.434 75.366 8.462 75.529 ;
      END
   END FE_OFN5889_n_41535

   PIN FE_OFN5896_n_143186
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.146 0.163 68.174 ;
      END
   END FE_OFN5896_n_143186

   PIN FE_OFN5963_n_41544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.05 0.163 64.078 ;
      END
   END FE_OFN5963_n_41544

   PIN FE_OFN9229_delay_add_ln34_unr2_unr4_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.402 75.366 76.43 75.529 ;
      END
   END FE_OFN9229_delay_add_ln34_unr2_unr4_stage2_stallmux_q_15_

   PIN FE_OFN9234_delay_add_ln34_unr2_unr2_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END FE_OFN9234_delay_add_ln34_unr2_unr2_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr6_unr0_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.626 75.366 8.654 75.529 ;
      END
   END delay_mul_ln34_unr6_unr0_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr6_unr3_stage2_stallmux_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.458 0.163 73.486 ;
      END
   END delay_mul_ln34_unr6_unr3_stage2_stallmux_z_3_

   PIN delay_mul_ln34_unr6_unr3_stage2_stallmux_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.466 75.366 4.494 75.529 ;
      END
   END delay_mul_ln34_unr6_unr3_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr6_unr3_stage2_stallmux_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.922 0.163 71.95 ;
      END
   END delay_mul_ln34_unr6_unr3_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr6_unr3_stage2_stallmux_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.538 0.163 71.566 ;
      END
   END delay_mul_ln34_unr6_unr3_stage2_stallmux_z_6_

   PIN delay_mul_ln34_unr6_unr3_stage2_stallmux_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.522 0.163 65.55 ;
      END
   END delay_mul_ln34_unr6_unr3_stage2_stallmux_z_7_

   PIN delay_mul_ln34_unr6_unr4_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 73.202 85.568 73.23 ;
      END
   END delay_mul_ln34_unr6_unr4_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr6_unr4_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 67.762 85.568 67.79 ;
      END
   END delay_mul_ln34_unr6_unr4_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr6_unr4_stage2_stallmux_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 44.786 85.568 44.814 ;
      END
   END delay_mul_ln34_unr6_unr4_stage2_stallmux_z_3_

   PIN mul_4685_72_n_127
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.602 0.163 71.63 ;
      END
   END mul_4685_72_n_127

   PIN mul_4685_72_n_153
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.922 0.163 55.95 ;
      END
   END mul_4685_72_n_153

   PIN mul_4685_72_n_81
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.738 75.366 2.766 75.529 ;
      END
   END mul_4685_72_n_81

   PIN mul_4685_72_n_848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.146 0.163 52.174 ;
      END
   END mul_4685_72_n_848

   PIN mul_4686_72_n_172
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.658 0.163 52.686 ;
      END
   END mul_4686_72_n_172

   PIN mul_4686_72_n_173
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.986 0.163 56.014 ;
      END
   END mul_4686_72_n_173

   PIN mul_4686_72_n_174
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.466 0.163 52.494 ;
      END
   END mul_4686_72_n_174

   PIN mul_4686_72_n_175
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.21 0.163 52.238 ;
      END
   END mul_4686_72_n_175

   PIN mul_4686_72_n_59
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.074 0.163 41.102 ;
      END
   END mul_4686_72_n_59

   PIN mul_4686_72_n_760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.138 0.163 41.166 ;
      END
   END mul_4686_72_n_760

   PIN mul_4686_72_n_765
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.946 0.163 40.974 ;
      END
   END mul_4686_72_n_765

   PIN mul_4686_72_n_825
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.818 0.163 40.846 ;
      END
   END mul_4686_72_n_825

   PIN mul_4692_72_n_100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.866 75.366 2.894 75.529 ;
      END
   END mul_4692_72_n_100

   PIN mul_4692_72_n_101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.738 75.366 2.766 75.529 ;
      END
   END mul_4692_72_n_101

   PIN mul_4692_72_n_125
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.138 0.163 73.166 ;
      END
   END mul_4692_72_n_125

   PIN mul_4692_72_n_128
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.426 0.163 69.454 ;
      END
   END mul_4692_72_n_128

   PIN mul_4692_72_n_99
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.69 0.163 72.718 ;
      END
   END mul_4692_72_n_99

   PIN n_100492
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.362 0.163 69.39 ;
      END
   END n_100492

   PIN n_101343
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.338 0.163 68.366 ;
      END
   END n_101343

   PIN n_103771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 71.282 0.163 71.31 ;
      END
   END n_103771

   PIN n_103826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.898 75.366 14.926 75.529 ;
      END
   END n_103826

   PIN n_104062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.37 0.163 48.398 ;
      END
   END n_104062

   PIN n_104069
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.658 0.163 44.686 ;
      END
   END n_104069

   PIN n_106541
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.722 0.163 44.75 ;
      END
   END n_106541

   PIN n_109205
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.866 75.366 10.894 75.529 ;
      END
   END n_109205

   PIN n_109222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.21 75.366 12.238 75.529 ;
      END
   END n_109222

   PIN n_109223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.274 75.366 12.302 75.529 ;
      END
   END n_109223

   PIN n_110029
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.674 75.366 18.702 75.529 ;
      END
   END n_110029

   PIN n_111074
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.762 75.366 19.79 75.529 ;
      END
   END n_111074

   PIN n_111156
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.754 0.163 72.782 ;
      END
   END n_111156

   PIN n_115715
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.53 0.163 52.558 ;
      END
   END n_115715

   PIN n_115716
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 52.466 0.163 52.494 ;
      END
   END n_115716

   PIN n_115759
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.37 0.163 56.398 ;
      END
   END n_115759

   PIN n_115760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.562 0.163 56.59 ;
      END
   END n_115760

   PIN n_115785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.402 0.163 60.43 ;
      END
   END n_115785

   PIN n_115786
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.626 0.163 56.654 ;
      END
   END n_115786

   PIN n_115911
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.89 0.163 59.918 ;
      END
   END n_115911

   PIN n_115923
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.434 0.163 48.462 ;
      END
   END n_115923

   PIN n_116134
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.786 0.163 44.814 ;
      END
   END n_116134

   PIN n_116475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.818 0.163 48.846 ;
      END
   END n_116475

   PIN n_116614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.602 0.163 63.63 ;
      END
   END n_116614

   PIN n_116752
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 56.306 0.163 56.334 ;
      END
   END n_116752

   PIN n_117032
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.626 0.163 48.654 ;
      END
   END n_117032

   PIN n_117103
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 44.658 0.163 44.686 ;
      END
   END n_117103

   PIN n_117106
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.802 75.366 2.83 75.529 ;
      END
   END n_117106

   PIN n_117107
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.802 75.366 2.83 75.529 ;
      END
   END n_117107

   PIN n_118624
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.954 0.163 59.982 ;
      END
   END n_118624

   PIN n_118625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.05 0.163 56.078 ;
      END
   END n_118625

   PIN n_118635
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.85 0.163 60.878 ;
      END
   END n_118635

   PIN n_118682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.498 0.163 48.526 ;
      END
   END n_118682

   PIN n_118902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.114 0.163 56.142 ;
      END
   END n_118902

   PIN n_118915
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.178 0.163 56.206 ;
      END
   END n_118915

   PIN n_119242
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 44.722 0.163 44.75 ;
      END
   END n_119242

   PIN n_119264
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.466 0.163 60.494 ;
      END
   END n_119264

   PIN n_119265
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.018 0.163 60.046 ;
      END
   END n_119265

   PIN n_119270
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.274 0.163 52.302 ;
      END
   END n_119270

   PIN n_120529
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 56.37 0.163 56.398 ;
      END
   END n_120529

   PIN n_121375
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.562 0.163 48.59 ;
      END
   END n_121375

   PIN n_122150
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 44.786 0.163 44.814 ;
      END
   END n_122150

   PIN n_122430
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.402 0.163 44.43 ;
      END
   END n_122430

   PIN n_123046
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.466 0.163 44.494 ;
      END
   END n_123046

   PIN n_123047
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.53 0.163 44.558 ;
      END
   END n_123047

   PIN n_123456
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 52.274 0.163 52.302 ;
      END
   END n_123456

   PIN n_127398
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.242 0.163 56.27 ;
      END
   END n_127398

   PIN n_127918
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 21.746 85.568 21.774 ;
      END
   END n_127918

   PIN n_128538
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.882 0.163 40.91 ;
      END
   END n_128538

   PIN n_128751
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.946 0.163 40.974 ;
      END
   END n_128751

   PIN n_129373
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 56.434 0.163 56.462 ;
      END
   END n_129373

   PIN n_130437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.338 0.163 52.366 ;
      END
   END n_130437

   PIN n_131022
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.882 0.163 40.91 ;
      END
   END n_131022

   PIN n_137688
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 72.562 85.568 72.59 ;
      END
   END n_137688

   PIN n_137761
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 56.242 85.568 56.27 ;
      END
   END n_137761

   PIN n_137849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.034 75.366 66.062 75.529 ;
      END
   END n_137849

   PIN n_35702
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.722 0.163 52.75 ;
      END
   END n_35702

   PIN n_36064
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.858 0.163 63.886 ;
      END
   END n_36064

   PIN n_37197
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 38.642 85.568 38.67 ;
      END
   END n_37197

   PIN n_37198
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.058 75.366 83.086 75.529 ;
      END
   END n_37198

   PIN n_37774
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 72.882 85.568 72.91 ;
      END
   END n_37774

   PIN n_37935
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.954 0.163 67.982 ;
      END
   END n_37935

   PIN n_37980
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 70.322 0.163 70.35 ;
      END
   END n_37980

   PIN n_38025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.082 0.163 60.11 ;
      END
   END n_38025

   PIN n_38471
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.018 0.163 68.046 ;
      END
   END n_38471

   PIN n_38472
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.082 0.163 68.11 ;
      END
   END n_38472

   PIN n_38617
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.002 0.163 70.03 ;
      END
   END n_38617

   PIN n_38618
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.066 0.163 70.094 ;
      END
   END n_38618

   PIN n_41119
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.25 75.366 3.278 75.529 ;
      END
   END n_41119

   PIN n_41226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.97 75.366 17.998 75.529 ;
      END
   END n_41226

   PIN n_41377
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 41.842 85.568 41.87 ;
      END
   END n_41377

   PIN n_43201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.778 75.366 17.806 75.529 ;
      END
   END n_43201

   PIN n_43202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.714 75.366 17.742 75.529 ;
      END
   END n_43202

   PIN n_43396
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.602 75.366 15.63 75.529 ;
      END
   END n_43396

   PIN n_43481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.61 75.366 18.638 75.529 ;
      END
   END n_43481

   PIN n_43848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.242 75.366 16.27 75.529 ;
      END
   END n_43848

   PIN n_44677
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.306 0.163 72.334 ;
      END
   END n_44677

   PIN n_44678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.234 75.366 21.262 75.529 ;
      END
   END n_44678

   PIN n_45925
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.05 0.163 72.078 ;
      END
   END n_45925

   PIN n_46856
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.914 0.163 60.942 ;
      END
   END n_46856

   PIN n_47058
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.922 0.163 63.95 ;
      END
   END n_47058

   PIN n_47110
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 67.826 0.163 67.854 ;
      END
   END n_47110

   PIN n_47630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.01 0.163 41.038 ;
      END
   END n_47630

   PIN n_47819
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.402 0.163 52.43 ;
      END
   END n_47819

   PIN n_50683
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.106 0.163 45.134 ;
      END
   END n_50683

   PIN n_50905
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.69 0.163 72.718 ;
      END
   END n_50905

   PIN n_51557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.498 0.163 72.526 ;
      END
   END n_51557

   PIN n_51614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 67.89 0.163 67.918 ;
      END
   END n_51614

   PIN n_52269
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 67.954 0.163 67.982 ;
      END
   END n_52269

   PIN n_52441
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.938 0.0 13.966 0.163 ;
      END
   END n_52441

   PIN n_52523
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.01 75.366 9.038 75.529 ;
      END
   END n_52523

   PIN n_53127
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.554 75.366 21.582 75.529 ;
      END
   END n_53127

   PIN n_53989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.626 0.163 48.654 ;
      END
   END n_53989

   PIN n_53990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.882 0.163 48.91 ;
      END
   END n_53990

   PIN n_53991
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.802 0.0 82.83 0.163 ;
      END
   END n_53991

   PIN n_54177
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.146 0.163 60.174 ;
      END
   END n_54177

   PIN n_55834
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.594 0.163 52.622 ;
      END
   END n_55834

   PIN n_56504
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.586 0.163 25.614 ;
      END
   END n_56504

   PIN n_56505
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.266 0.163 33.294 ;
      END
   END n_56505

   PIN n_57641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.682 75.366 21.71 75.529 ;
      END
   END n_57641

   PIN n_58613
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.69 0.163 48.718 ;
      END
   END n_58613

   PIN n_58614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 65.266 0.163 65.294 ;
      END
   END n_58614

   PIN n_58621
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.21 0.163 60.238 ;
      END
   END n_58621

   PIN n_58622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.306 0.163 64.334 ;
      END
   END n_58622

   PIN n_62348
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.434 0.163 56.462 ;
      END
   END n_62348

   PIN n_62349
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.986 0.163 64.014 ;
      END
   END n_62349

   PIN n_63582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.85 0.163 44.878 ;
      END
   END n_63582

   PIN n_64651
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.914 0.163 44.942 ;
      END
   END n_64651

   PIN n_65851
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 52.338 0.163 52.366 ;
      END
   END n_65851

   PIN n_76609
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 44.85 0.163 44.878 ;
      END
   END n_76609

   PIN n_84147
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.066 75.366 22.094 75.529 ;
      END
   END n_84147

   PIN n_88793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.306 0.163 56.334 ;
      END
   END n_88793

   PIN n_89861
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.298 75.366 21.326 75.529 ;
      END
   END n_89861

   PIN n_90532
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.41 75.366 23.438 75.529 ;
      END
   END n_90532

   PIN n_94236
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.154 75.366 15.182 75.529 ;
      END
   END n_94236

   PIN n_96014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.434 0.163 72.462 ;
      END
   END n_96014

   PIN n_96031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.242 0.163 72.27 ;
      END
   END n_96031

   PIN n_96563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.69 0.163 48.718 ;
      END
   END n_96563

   PIN n_98744
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.978 0.163 45.006 ;
      END
   END n_98744

   PIN n_98745
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.042 0.163 45.07 ;
      END
   END n_98745

   PIN FE_OCPN15689_FE_OFN12113_n_41363
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.794 0.163 63.822 ;
      END
   END FE_OCPN15689_FE_OFN12113_n_41363

   PIN FE_OFN1071_n_16034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.122 0.0 83.15 0.163 ;
      END
   END FE_OFN1071_n_16034

   PIN FE_OFN11840_n_144163
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.882 75.447 8.91 75.529 ;
      END
   END FE_OFN11840_n_144163

   PIN FE_OFN11843_n_144163
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.634 75.447 19.662 75.529 ;
      END
   END FE_OFN11843_n_144163

   PIN FE_OFN11845_n_144163
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.922 75.366 23.95 75.529 ;
      END
   END FE_OFN11845_n_144163

   PIN FE_OFN11848_n_144163
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.794 0.082 63.822 ;
      END
   END FE_OFN11848_n_144163

   PIN FE_OFN12052_n_41878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.794 75.366 23.822 75.529 ;
      END
   END FE_OFN12052_n_41878

   PIN FE_OFN12068_n_41544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.154 75.366 23.182 75.529 ;
      END
   END FE_OFN12068_n_41544

   PIN FE_OFN12094_n_41679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.218 75.366 15.246 75.529 ;
      END
   END FE_OFN12094_n_41679

   PIN FE_OFN12111_n_41363
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.098 75.366 18.126 75.529 ;
      END
   END FE_OFN12111_n_41363

   PIN FE_OFN12995_n_41504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.402 75.447 4.43 75.529 ;
      END
   END FE_OFN12995_n_41504

   PIN FE_OFN13259_n_143327
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.234 75.366 13.262 75.529 ;
      END
   END FE_OFN13259_n_143327

   PIN FE_OFN13274_n_143160
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.178 75.366 24.206 75.529 ;
      END
   END FE_OFN13274_n_143160

   PIN FE_OFN13276_n_143160
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.73 0.163 63.758 ;
      END
   END FE_OFN13276_n_143160

   PIN FE_OFN13280_n_143159
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.234 75.366 29.262 75.529 ;
      END
   END FE_OFN13280_n_143159

   PIN FE_OFN13679_n_143468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.962 75.366 22.99 75.529 ;
      END
   END FE_OFN13679_n_143468

   PIN FE_OFN13684_n_143467
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.818 75.366 16.846 75.529 ;
      END
   END FE_OFN13684_n_143467

   PIN FE_OFN13697_n_143411
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.594 75.447 12.622 75.529 ;
      END
   END FE_OFN13697_n_143411

   PIN FE_OFN13720_n_143132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.41 0.082 71.438 ;
      END
   END FE_OFN13720_n_143132

   PIN FE_OFN13725_n_143131
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.266 75.366 25.294 75.529 ;
      END
   END FE_OFN13725_n_143131

   PIN FE_OFN13770_n_41154
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.01 75.366 9.038 75.529 ;
      END
   END FE_OFN13770_n_41154

   PIN FE_OFN13784_n_41769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.786 0.163 52.814 ;
      END
   END FE_OFN13784_n_41769

   PIN FE_OFN13836_n_143217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.53 0.163 60.558 ;
      END
   END FE_OFN13836_n_143217

   PIN FE_OFN13840_n_143189
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.37 0.163 64.398 ;
      END
   END FE_OFN13840_n_143189

   PIN FE_OFN13920_n_143215
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.074 75.366 9.102 75.529 ;
      END
   END FE_OFN13920_n_143215

   PIN FE_OFN13926_n_143214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.234 75.366 5.262 75.529 ;
      END
   END FE_OFN13926_n_143214

   PIN FE_OFN13933_n_143213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.178 0.163 64.206 ;
      END
   END FE_OFN13933_n_143213

   PIN FE_OFN13937_n_143187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.93 75.366 2.958 75.529 ;
      END
   END FE_OFN13937_n_143187

   PIN FE_OFN13942_n_143186
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.562 0.163 48.59 ;
      END
   END FE_OFN13942_n_143186

   PIN FE_OFN13948_n_143185
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.498 75.366 32.526 75.529 ;
      END
   END FE_OFN13948_n_143185

   PIN FE_OFN13949_n_143185
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.858 0.163 55.886 ;
      END
   END FE_OFN13949_n_143185

   PIN FE_OFN13970_n_41362
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.042 75.366 21.07 75.529 ;
      END
   END FE_OFN13970_n_41362

   PIN FE_OFN13979_n_41537
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.474 75.366 7.502 75.529 ;
      END
   END FE_OFN13979_n_41537

   PIN FE_OFN14343_n_67347
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.218 75.366 23.246 75.529 ;
      END
   END FE_OFN14343_n_67347

   PIN FE_OFN14412_n_41429
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.786 75.366 20.814 75.529 ;
      END
   END FE_OFN14412_n_41429

   PIN FE_OFN14553_n_67346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.682 75.366 21.71 75.529 ;
      END
   END FE_OFN14553_n_67346

   PIN FE_OFN15019_n_41544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.93 75.366 2.958 75.529 ;
      END
   END FE_OFN15019_n_41544

   PIN FE_OFN15033_n_41535
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.882 75.366 16.91 75.529 ;
      END
   END FE_OFN15033_n_41535

   PIN FE_OFN15038_n_41507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.162 75.366 10.19 75.529 ;
      END
   END FE_OFN15038_n_41507

   PIN FE_OFN15281_n_67352
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.146 0.163 68.174 ;
      END
   END FE_OFN15281_n_67352

   PIN FE_OFN16051_n_67347
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 69.746 0.163 69.774 ;
      END
   END FE_OFN16051_n_67347

   PIN FE_OFN4352_n_67017
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.914 0.0 4.942 0.163 ;
      END
   END FE_OFN4352_n_67017

   PIN FE_OFN5763_n_41506
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.826 75.366 19.854 75.529 ;
      END
   END FE_OFN5763_n_41506

   PIN FE_OFN5823_n_143157
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.026 75.366 31.054 75.529 ;
      END
   END FE_OFN5823_n_143157

   PIN FE_OFN5854_n_143129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.138 75.366 9.166 75.529 ;
      END
   END FE_OFN5854_n_143129

   PIN FE_OFN5871_n_143132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.25 75.366 19.278 75.529 ;
      END
   END FE_OFN5871_n_143132

   PIN FE_OFN5873_n_41152
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.754 75.447 8.782 75.529 ;
      END
   END FE_OFN5873_n_41152

   PIN FE_OFN5877_n_143130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.074 75.366 33.102 75.529 ;
      END
   END FE_OFN5877_n_143130

   PIN FE_OFN5908_n_41536
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.97 75.366 9.998 75.529 ;
      END
   END FE_OFN5908_n_41536

   PIN FE_OFN5950_n_41543
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.346 75.366 15.374 75.529 ;
      END
   END FE_OFN5950_n_41543

   PIN FE_OFN5982_n_143325
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.426 75.447 29.454 75.529 ;
      END
   END FE_OFN5982_n_143325

   PIN FE_OFN6009_n_41879
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.274 0.163 68.302 ;
      END
   END FE_OFN6009_n_41879

   PIN FE_OFN6021_n_41878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.098 75.366 26.126 75.529 ;
      END
   END FE_OFN6021_n_41878

   PIN FE_OFN6057_n_140218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.21 75.366 20.238 75.529 ;
      END
   END FE_OFN6057_n_140218

   PIN FE_OFN6076_n_67348
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.594 0.163 68.622 ;
      END
   END FE_OFN6076_n_67348

   PIN FE_OFN6139_n_67344
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.186 75.366 19.214 75.529 ;
      END
   END FE_OFN6139_n_67344

   PIN FE_OFN9228_delay_add_ln34_unr2_unr4_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.722 0.163 36.75 ;
      END
   END FE_OFN9228_delay_add_ln34_unr2_unr4_stage2_stallmux_q_15_

   PIN b_6_1_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.186 75.447 3.214 75.529 ;
      END
   END b_6_1_5

   PIN b_6_1_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.122 75.366 3.15 75.529 ;
      END
   END b_6_1_6

   PIN b_6_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.338 0.082 68.366 ;
      END
   END b_6_3_0

   PIN b_6_3_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.554 0.082 69.582 ;
      END
   END b_6_3_1

   PIN b_6_3_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.338 0.163 60.366 ;
      END
   END b_6_3_2

   PIN b_6_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.498 75.447 8.526 75.529 ;
      END
   END b_6_3_3

   PIN b_6_3_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.994 75.366 3.022 75.529 ;
      END
   END b_6_3_5

   PIN b_6_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.866 0.0 34.894 0.082 ;
      END
   END b_6_4_0

   PIN b_6_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.354 75.447 34.382 75.529 ;
      END
   END b_6_4_1

   PIN b_6_4_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.266 75.366 17.294 75.529 ;
      END
   END b_6_4_10

   PIN b_6_4_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.298 75.366 29.326 75.529 ;
      END
   END b_6_4_12

   PIN b_6_4_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.538 75.447 31.566 75.529 ;
      END
   END b_6_4_2

   PIN b_6_4_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.53 75.447 28.558 75.529 ;
      END
   END b_6_4_3

   PIN b_6_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 65.522 0.082 65.55 ;
      END
   END b_6_4_4

   PIN b_6_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 67.634 0.082 67.662 ;
      END
   END b_6_4_5

   PIN b_6_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.69 0.163 56.718 ;
      END
   END b_6_4_6

   PIN b_6_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.706 75.366 30.734 75.529 ;
      END
   END b_6_4_7

   PIN b_6_4_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.898 0.0 30.926 0.163 ;
      END
   END b_6_4_8

   PIN b_6_4_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.242 0.163 64.27 ;
      END
   END b_6_4_9

   PIN b_6_8_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.314 75.366 19.342 75.529 ;
      END
   END b_6_8_0

   PIN b_6_8_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.666 75.366 15.694 75.529 ;
      END
   END b_6_8_10

   PIN b_6_8_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.378 75.366 19.406 75.529 ;
      END
   END b_6_8_11

   PIN b_6_8_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.89 75.366 19.918 75.529 ;
      END
   END b_6_8_13

   PIN b_6_8_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.346 75.366 23.374 75.529 ;
      END
   END b_6_8_2

   PIN b_6_8_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.442 75.366 19.47 75.529 ;
      END
   END b_6_8_3

   PIN b_6_8_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.762 75.366 19.79 75.529 ;
      END
   END b_6_8_4

   PIN b_6_8_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.298 75.366 21.326 75.529 ;
      END
   END b_6_8_5

   PIN b_6_8_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.946 75.366 16.974 75.529 ;
      END
   END b_6_8_6

   PIN b_6_8_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.474 75.366 15.502 75.529 ;
      END
   END b_6_8_7

   PIN b_6_8_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.282 75.366 15.31 75.529 ;
      END
   END b_6_8_8

   PIN b_6_8_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.114 75.366 16.142 75.529 ;
      END
   END b_6_8_9

   PIN delay_add_ln34_unr2_unr2_stage2_stallmux_q_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 0.946 85.568 0.974 ;
      END
   END delay_add_ln34_unr2_unr2_stage2_stallmux_q_13_

   PIN delay_add_ln34_unr2_unr2_stage2_stallmux_q_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 16.242 85.568 16.27 ;
      END
   END delay_add_ln34_unr2_unr2_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr6_unr0_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.922 75.366 7.95 75.529 ;
      END
   END delay_mul_ln34_unr6_unr0_stage2_stallmux_z_7_

   PIN delay_mul_ln34_unr6_unr8_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.29 75.366 42.318 75.529 ;
      END
   END delay_mul_ln34_unr6_unr8_stage2_stallmux_z_2_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.954 75.447 43.982 75.529 ;
      END
   END ispd_clk

   PIN mul_4384_72_n_322
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 47.602 85.568 47.63 ;
      END
   END mul_4384_72_n_322

   PIN mul_4385_72_n_291
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.186 0.0 83.214 0.163 ;
      END
   END mul_4385_72_n_291

   PIN mul_4385_72_n_293
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 37.362 85.568 37.39 ;
      END
   END mul_4385_72_n_293

   PIN mul_4685_72_n_113
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.394 0.163 73.422 ;
      END
   END mul_4685_72_n_113

   PIN mul_4685_72_n_114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.826 75.366 3.854 75.529 ;
      END
   END mul_4685_72_n_114

   PIN mul_4685_72_n_123
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.01 0.163 73.038 ;
      END
   END mul_4685_72_n_123

   PIN mul_4685_72_n_124
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.754 0.163 72.782 ;
      END
   END mul_4685_72_n_124

   PIN mul_4685_72_n_126
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.282 0.163 71.31 ;
      END
   END mul_4685_72_n_126

   PIN mul_4685_72_n_128
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.45 0.163 70.478 ;
      END
   END mul_4685_72_n_128

   PIN mul_4686_72_n_75
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.754 0.163 40.782 ;
      END
   END mul_4686_72_n_75

   PIN n_100517
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.002 75.366 14.03 75.529 ;
      END
   END n_100517

   PIN n_100894
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.666 0.163 63.694 ;
      END
   END n_100894

   PIN n_100908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 65.33 0.163 65.358 ;
      END
   END n_100908

   PIN n_103167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.538 0.163 63.566 ;
      END
   END n_103167

   PIN n_104067
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.114 0.163 64.142 ;
      END
   END n_104067

   PIN n_104070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.594 0.163 44.622 ;
      END
   END n_104070

   PIN n_105146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.178 0.163 72.206 ;
      END
   END n_105146

   PIN n_107966
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 61.042 0.163 61.07 ;
      END
   END n_107966

   PIN n_109265
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.506 75.366 27.534 75.529 ;
      END
   END n_109265

   PIN n_110663
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.37 0.163 72.398 ;
      END
   END n_110663

   PIN n_110915
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.562 75.366 16.59 75.529 ;
      END
   END n_110915

   PIN n_112026
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.33 0.163 73.358 ;
      END
   END n_112026

   PIN n_116135
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.306 0.163 48.334 ;
      END
   END n_116135

   PIN n_116476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.498 0.163 48.526 ;
      END
   END n_116476

   PIN n_122251
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 55.282 85.568 55.31 ;
      END
   END n_122251

   PIN n_123110
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.602 0.163 63.63 ;
      END
   END n_123110

   PIN n_123111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.826 0.163 59.854 ;
      END
   END n_123111

   PIN n_125285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 55.346 85.568 55.374 ;
      END
   END n_125285

   PIN n_125286
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.122 75.366 83.15 75.529 ;
      END
   END n_125286

   PIN n_126760
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.754 0.163 48.782 ;
      END
   END n_126760

   PIN n_140296
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 85.405 6.322 85.568 6.35 ;
      END
   END n_140296

   PIN n_143329
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.514 75.447 6.542 75.529 ;
      END
   END n_143329

   PIN n_143413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.13 75.447 6.158 75.529 ;
      END
   END n_143413

   PIN n_143595
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 67.762 0.163 67.79 ;
      END
   END n_143595

   PIN n_143865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.978 0.163 61.006 ;
      END
   END n_143865

   PIN n_31805
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.266 0.163 73.294 ;
      END
   END n_31805

   PIN n_33135
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.426 0.163 29.454 ;
      END
   END n_33135

   PIN n_34106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.058 75.366 3.086 75.529 ;
      END
   END n_34106

   PIN n_34265
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.106 0.163 37.134 ;
      END
   END n_34265

   PIN n_34503
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.378 75.366 3.406 75.529 ;
      END
   END n_34503

   PIN n_34853
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.866 75.366 2.894 75.529 ;
      END
   END n_34853

   PIN n_35129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.746 0.163 21.774 ;
      END
   END n_35129

   PIN n_35323
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.042 0.163 37.07 ;
      END
   END n_35323

   PIN n_36377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.25 75.366 83.278 75.529 ;
      END
   END n_36377

   PIN n_37528
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.818 0.163 72.846 ;
      END
   END n_37528

   PIN n_37611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.202 0.163 73.23 ;
      END
   END n_37611

   PIN n_37704
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.21 0.163 68.238 ;
      END
   END n_37704

   PIN n_38380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.082 0.163 68.11 ;
      END
   END n_38380

   PIN n_41039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.474 0.163 63.502 ;
      END
   END n_41039

   PIN n_41241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.146 75.366 20.174 75.529 ;
      END
   END n_41241

   PIN n_41333
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.882 0.163 72.91 ;
      END
   END n_41333

   PIN n_41505
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.522 75.366 9.55 75.529 ;
      END
   END n_41505

   PIN n_41698
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.722 75.366 20.75 75.529 ;
      END
   END n_41698

   PIN n_43847
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.538 75.366 15.566 75.529 ;
      END
   END n_43847

   PIN n_44259
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.834 75.366 22.862 75.529 ;
      END
   END n_44259

   PIN n_46640
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.33 75.366 17.358 75.529 ;
      END
   END n_46640

   PIN n_47006
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.89 0.163 67.918 ;
      END
   END n_47006

   PIN n_47088
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.786 0.163 60.814 ;
      END
   END n_47088

   PIN n_47111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.826 0.163 67.854 ;
      END
   END n_47111

   PIN n_47947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.498 0.163 56.526 ;
      END
   END n_47947

   PIN n_49044
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.426 75.366 21.454 75.529 ;
      END
   END n_49044

   PIN n_49385
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.698 75.366 3.726 75.529 ;
      END
   END n_49385

   PIN n_52268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.538 0.163 63.566 ;
      END
   END n_52268

   PIN n_52442
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.482 0.163 2.51 ;
      END
   END n_52442

   PIN n_52806
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.666 75.366 23.694 75.529 ;
      END
   END n_52806

   PIN n_53026
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.274 0.163 60.302 ;
      END
   END n_53026

   PIN n_53126
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.618 75.366 21.646 75.529 ;
      END
   END n_53126

   PIN n_55075
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.818 0.163 72.846 ;
      END
   END n_55075

   PIN n_55277
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.794 75.366 15.822 75.529 ;
      END
   END n_55277

   PIN n_55441
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.834 75.366 14.862 75.529 ;
      END
   END n_55441

   PIN n_56027
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 66.802 0.163 66.83 ;
      END
   END n_56027

   PIN n_57044
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.746 75.366 21.774 75.529 ;
      END
   END n_57044

   PIN n_57047
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.554 75.366 21.582 75.529 ;
      END
   END n_57047

   PIN n_58615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 67.122 0.163 67.15 ;
      END
   END n_58615

   PIN n_76128
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 68.018 0.163 68.046 ;
      END
   END n_76128

   PIN n_80052
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.626 75.366 16.654 75.529 ;
      END
   END n_80052

   PIN n_80708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.082 0.163 52.11 ;
      END
   END n_80708

   PIN n_81744
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.434 75.366 16.462 75.529 ;
      END
   END n_81744

   PIN n_82461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.762 0.163 59.79 ;
      END
   END n_82461

   PIN n_83267
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.17 75.366 13.198 75.529 ;
      END
   END n_83267

   PIN n_85057
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.306 75.366 16.334 75.529 ;
      END
   END n_85057

   PIN n_89837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.762 0.163 67.79 ;
      END
   END n_89837

   PIN n_89839
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.026 75.366 15.054 75.529 ;
      END
   END n_89839

   PIN n_90520
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.666 0.163 63.694 ;
      END
   END n_90520

   PIN n_90524
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 52.402 0.163 52.43 ;
      END
   END n_90524

   PIN n_92013
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.426 75.366 13.454 75.529 ;
      END
   END n_92013

   PIN n_94239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.066 75.366 22.094 75.529 ;
      END
   END n_94239

   PIN n_94241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.002 75.366 22.03 75.529 ;
      END
   END n_94241

   PIN n_96030
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.042 75.366 13.07 75.529 ;
      END
   END n_96030

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 85.568 75.53 ;
      LAYER V1 ;
         RECT 0.0 0.0 85.568 75.53 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 85.568 75.53 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 85.568 75.53 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 85.568 75.53 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 85.568 75.53 ;
      LAYER M1 ;
         RECT 0.0 0.0 85.568 75.53 ;
   END
END h9_mgc_matrix_mult_b

MACRO h8_mgc_matrix_mult_b
   CLASS BLOCK ;
   FOREIGN h8 ;
   ORIGIN 0 0 ;
   SIZE 99.456 BY 107.52 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN15134_n_30145
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 52.466 0.163 52.494 ;
      END
   END FE_OFN15134_n_30145

   PIN FE_OFN15136_n_31158
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 88.562 0.163 88.59 ;
      END
   END FE_OFN15136_n_31158

   PIN FE_OFN16292_n_22751
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.074 0.0 33.102 0.163 ;
      END
   END FE_OFN16292_n_22751

   PIN FE_OFN17812_delay_mul_ln34_unr7_unr9_stage2_stallmux_z_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.914 0.0 12.942 0.163 ;
      END
   END FE_OFN17812_delay_mul_ln34_unr7_unr9_stage2_stallmux_z_11_

   PIN FE_OFN17822_n_137819
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.69 0.0 40.718 0.163 ;
      END
   END FE_OFN17822_n_137819

   PIN FE_OFN18396_n_31131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.778 107.357 17.806 107.52 ;
      END
   END FE_OFN18396_n_31131

   PIN FE_OFN18402_n_30571
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.442 107.357 19.47 107.52 ;
      END
   END FE_OFN18402_n_30571

   PIN FE_OFN18458_n_29943
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.626 107.357 0.654 107.52 ;
      END
   END FE_OFN18458_n_29943

   PIN FE_OFN18462_n_28644
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.762 0.163 59.79 ;
      END
   END FE_OFN18462_n_28644

   PIN FE_OFN18464_n_28105
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.202 0.163 57.23 ;
      END
   END FE_OFN18464_n_28105

   PIN FE_OFN18466_n_27225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 54.002 0.163 54.03 ;
      END
   END FE_OFN18466_n_27225

   PIN FE_OFN6270_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.914 0.0 36.942 0.163 ;
      END
   END FE_OFN6270_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_10_

   PIN FE_OFN6274_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.538 0.0 71.566 0.163 ;
      END
   END FE_OFN6274_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_9_

   PIN FE_OFN6330_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.602 0.0 71.63 0.163 ;
      END
   END FE_OFN6330_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_8_

   PIN FE_OFN6338_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.162 0.0 42.19 0.163 ;
      END
   END FE_OFN6338_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_6_

   PIN FE_OFN6340_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.602 0.0 71.63 0.163 ;
      END
   END FE_OFN6340_delay_mul_ln34_unr7_unr4_stage2_stallmux_z_5_

   PIN FE_OFN8209_n_30818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.546 0.163 98.574 ;
      END
   END FE_OFN8209_n_30818

   PIN FE_OFN8218_n_31243
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.178 107.357 40.206 107.52 ;
      END
   END FE_OFN8218_n_31243

   PIN FE_OFN8458_n_27222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 81.522 0.163 81.55 ;
      END
   END FE_OFN8458_n_27222

   PIN FE_OFN8463_n_25371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.962 0.163 62.99 ;
      END
   END FE_OFN8463_n_25371

   PIN FE_OFN8467_n_24044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.898 0.163 86.926 ;
      END
   END FE_OFN8467_n_24044

   PIN FE_OFN8627_n_30345
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.298 107.357 37.326 107.52 ;
      END
   END FE_OFN8627_n_30345

   PIN FE_OFN8630_n_30620
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.322 0.163 94.35 ;
      END
   END FE_OFN8630_n_30620

   PIN FE_OFN8631_n_30852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.738 107.357 10.766 107.52 ;
      END
   END FE_OFN8631_n_30852

   PIN FE_OFN8633_n_31042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.042 0.163 77.07 ;
      END
   END FE_OFN8633_n_31042

   PIN FE_OFN8640_n_30028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.402 107.357 36.43 107.52 ;
      END
   END FE_OFN8640_n_30028

   PIN FE_OFN8642_n_29615
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.642 0.163 94.67 ;
      END
   END FE_OFN8642_n_29615

   PIN FE_OFN8663_n_28865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.522 0.163 25.55 ;
      END
   END FE_OFN8663_n_28865

   PIN FE_OFN8665_n_29329
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.682 0.163 21.71 ;
      END
   END FE_OFN8665_n_29329

   PIN FE_OFN8668_n_30136
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.642 0.0 38.67 0.163 ;
      END
   END FE_OFN8668_n_30136

   PIN FE_OFN8673_n_27200
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.138 0.0 33.166 0.163 ;
      END
   END FE_OFN8673_n_27200

   PIN FE_OFN8689_n_6646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.426 0.0 29.454 0.163 ;
      END
   END FE_OFN8689_n_6646

   PIN FE_OFN8711_n_27536
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.482 0.163 58.51 ;
      END
   END FE_OFN8711_n_27536

   PIN FE_OFN8834_n_25354
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.594 0.0 44.622 0.163 ;
      END
   END FE_OFN8834_n_25354

   PIN FE_OFN8838_n_24020
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.274 0.0 52.302 0.163 ;
      END
   END FE_OFN8838_n_24020

   PIN FE_OFN8841_n_22184
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.202 0.0 33.23 0.163 ;
      END
   END FE_OFN8841_n_22184

   PIN FE_OFN9032_n_18065
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.482 0.0 2.51 0.163 ;
      END
   END FE_OFN9032_n_18065

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.658 0.0 44.686 0.163 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_10_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.402 0.0 52.43 0.163 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_11_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.178 0.0 56.206 0.163 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.082 0.0 60.11 0.163 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.962 0.0 22.99 0.163 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.65 0.0 17.678 0.163 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.714 0.0 17.742 0.163 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_9_

   PIN delay_mul_ln34_unr7_unr2_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.362 0.0 29.39 0.163 ;
      END
   END delay_mul_ln34_unr7_unr2_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.378 0.0 75.406 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.642 0.0 94.67 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_11_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 83.122 0.0 83.15 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 28.402 99.456 28.43 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 30.322 99.456 30.35 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.93 0.0 90.958 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.666 0.0 71.694 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.442 0.0 75.47 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.442 0.0 75.47 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_3_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.962 0.0 86.99 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.706 0.0 94.734 0.163 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.242 0.0 56.27 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_10_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.242 0.0 56.27 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_11_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.826 0.0 35.854 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.626 0.0 48.654 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.922 0.0 63.95 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.722 0.0 44.75 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.29 0.0 10.318 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.402 0.0 52.43 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.362 0.0 29.39 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.306 0.0 56.334 0.163 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_q_9_

   PIN delay_mul_ln34_unr7_unr9_stage2_stallmux_z_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.322 0.0 6.35 0.163 ;
      END
   END delay_mul_ln34_unr7_unr9_stage2_stallmux_z_10_

   PIN delay_mul_ln34_unr7_unr9_stage2_stallmux_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.85 0.0 4.878 0.163 ;
      END
   END delay_mul_ln34_unr7_unr9_stage2_stallmux_z_6_

   PIN delay_mul_ln34_unr7_unr9_stage2_stallmux_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.17 0.0 5.198 0.163 ;
      END
   END delay_mul_ln34_unr7_unr9_stage2_stallmux_z_7_

   PIN delay_mul_ln34_unr7_unr9_stage2_stallmux_z_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 4.722 99.456 4.75 ;
      END
   END delay_mul_ln34_unr7_unr9_stage2_stallmux_z_8_

   PIN delay_mul_ln34_unr7_unr9_stage2_stallmux_z_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.722 0.0 4.75 0.163 ;
      END
   END delay_mul_ln34_unr7_unr9_stage2_stallmux_z_9_

   PIN delay_mul_ln34_unr8_unr7_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.866 0.163 18.894 ;
      END
   END delay_mul_ln34_unr8_unr7_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr9_unr6_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.378 0.0 35.406 0.163 ;
      END
   END delay_mul_ln34_unr9_unr6_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr9_unr6_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.306 0.0 32.334 0.163 ;
      END
   END delay_mul_ln34_unr9_unr6_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr9_unr6_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.754 0.0 32.782 0.163 ;
      END
   END delay_mul_ln34_unr9_unr6_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr9_unr6_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.658 0.0 20.686 0.163 ;
      END
   END delay_mul_ln34_unr9_unr6_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr9_unr6_stage2_stallmux_z_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.498 0.0 24.526 0.163 ;
      END
   END delay_mul_ln34_unr9_unr6_stage2_stallmux_z_10_

   PIN delay_mul_ln34_unr9_unr6_stage2_stallmux_z_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.226 0.0 42.254 0.163 ;
      END
   END delay_mul_ln34_unr9_unr6_stage2_stallmux_z_11_

   PIN delay_mul_ln34_unr9_unr6_stage2_stallmux_z_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.65 0.0 25.678 0.163 ;
      END
   END delay_mul_ln34_unr9_unr6_stage2_stallmux_z_9_

   PIN n_104375
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.938 0.163 13.966 ;
      END
   END n_104375

   PIN n_106153
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.066 0.163 14.094 ;
      END
   END n_106153

   PIN n_107402
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 84.082 0.163 84.11 ;
      END
   END n_107402

   PIN n_110538
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.578 0.163 6.606 ;
      END
   END n_110538

   PIN n_122192
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.666 0.163 79.694 ;
      END
   END n_122192

   PIN n_144102
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.138 0.0 25.166 0.163 ;
      END
   END n_144102

   PIN n_18141
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.786 0.0 44.814 0.163 ;
      END
   END n_18141

   PIN n_18874
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.842 107.357 17.87 107.52 ;
      END
   END n_18874

   PIN n_19306
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.218 0.0 15.246 0.163 ;
      END
   END n_19306

   PIN n_19638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.466 0.163 44.494 ;
      END
   END n_19638

   PIN n_19982
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.906 0.163 73.934 ;
      END
   END n_19982

   PIN n_19998
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 71.602 0.163 71.63 ;
      END
   END n_19998

   PIN n_21907
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.994 0.0 27.022 0.163 ;
      END
   END n_21907

   PIN n_23034
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.626 107.357 32.654 107.52 ;
      END
   END n_23034

   PIN n_23348
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.466 0.0 52.494 0.163 ;
      END
   END n_23348

   PIN n_23375
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.706 0.163 94.734 ;
      END
   END n_23375

   PIN n_24065
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.234 0.0 13.262 0.163 ;
      END
   END n_24065

   PIN n_24315
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.186 0.163 43.214 ;
      END
   END n_24315

   PIN n_24449
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.162 0.0 50.19 0.163 ;
      END
   END n_24449

   PIN n_24653
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.602 0.0 47.63 0.163 ;
      END
   END n_24653

   PIN n_24674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.282 0.163 79.31 ;
      END
   END n_24674

   PIN n_24729
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.418 0.0 50.446 0.163 ;
      END
   END n_24729

   PIN n_24782
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.906 0.0 49.934 0.163 ;
      END
   END n_24782

   PIN n_24783
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.778 0.0 49.806 0.163 ;
      END
   END n_24783

   PIN n_25168
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.05 0.0 48.078 0.163 ;
      END
   END n_25168

   PIN n_25376
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.282 0.163 39.31 ;
      END
   END n_25376

   PIN n_25386
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.338 0.0 12.366 0.163 ;
      END
   END n_25386

   PIN n_25409
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.61 0.163 98.638 ;
      END
   END n_25409

   PIN n_25453
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.642 0.0 94.67 0.163 ;
      END
   END n_25453

   PIN n_25807
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.178 0.0 48.206 0.163 ;
      END
   END n_25807

   PIN n_26004
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.178 107.357 80.206 107.52 ;
      END
   END n_26004

   PIN n_26006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.042 0.163 45.07 ;
      END
   END n_26006

   PIN n_26016
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.882 0.0 32.91 0.163 ;
      END
   END n_26016

   PIN n_26061
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.722 0.0 44.75 0.163 ;
      END
   END n_26061

   PIN n_26618
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.226 0.0 42.254 0.163 ;
      END
   END n_26618

   PIN n_26619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.658 0.0 44.686 0.163 ;
      END
   END n_26619

   PIN n_26638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 46.322 0.163 46.35 ;
      END
   END n_26638

   PIN n_26650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.386 0.163 102.414 ;
      END
   END n_26650

   PIN n_26651
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.946 0.0 32.974 0.163 ;
      END
   END n_26651

   PIN n_26674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.05 0.163 56.078 ;
      END
   END n_26674

   PIN n_27195
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.498 0.0 40.526 0.163 ;
      END
   END n_27195

   PIN n_27239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.154 0.0 15.182 0.163 ;
      END
   END n_27239

   PIN n_27295
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.146 0.163 60.174 ;
      END
   END n_27295

   PIN n_27323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.634 0.0 43.662 0.163 ;
      END
   END n_27323

   PIN n_27563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.01 0.0 33.038 0.163 ;
      END
   END n_27563

   PIN n_27656
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.626 0.0 24.654 0.163 ;
      END
   END n_27656

   PIN n_27657
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.69 0.0 24.718 0.163 ;
      END
   END n_27657

   PIN n_27696
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.242 0.0 40.27 0.163 ;
      END
   END n_27696

   PIN n_27719
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.754 0.0 40.782 0.163 ;
      END
   END n_27719

   PIN n_27864
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.45 0.163 102.478 ;
      END
   END n_27864

   PIN n_27896
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.882 0.163 48.91 ;
      END
   END n_27896

   PIN n_27914
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.906 0.0 41.934 0.163 ;
      END
   END n_27914

   PIN n_27936
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.114 0.0 40.142 0.163 ;
      END
   END n_27936

   PIN n_28388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.514 0.163 102.542 ;
      END
   END n_28388

   PIN n_28444
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.73 0.163 47.758 ;
      END
   END n_28444

   PIN n_28624
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.762 0.163 43.79 ;
      END
   END n_28624

   PIN n_28690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.322 0.163 46.35 ;
      END
   END n_28690

   PIN n_28758
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.402 0.163 44.43 ;
      END
   END n_28758

   PIN n_28891
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.322 107.357 6.35 107.52 ;
      END
   END n_28891

   PIN n_29119
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 0.754 107.357 0.782 107.52 ;
      END
   END n_29119

   PIN n_29177
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.338 0.163 52.366 ;
      END
   END n_29177

   PIN n_29352
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.674 0.163 98.702 ;
      END
   END n_29352

   PIN n_29433
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.338 0.0 36.366 0.163 ;
      END
   END n_29433

   PIN n_29550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.266 0.163 57.294 ;
      END
   END n_29550

   PIN n_29572
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.45 107.357 22.478 107.52 ;
      END
   END n_29572

   PIN n_29666
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.658 0.0 36.686 0.163 ;
      END
   END n_29666

   PIN n_29667
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.402 0.0 36.43 0.163 ;
      END
   END n_29667

   PIN n_29966
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.706 107.357 22.734 107.52 ;
      END
   END n_29966

   PIN n_30272
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.322 0.163 62.35 ;
      END
   END n_30272

   PIN n_30290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.21 107.357 20.238 107.52 ;
      END
   END n_30290

   PIN n_30440
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 3.442 99.456 3.47 ;
      END
   END n_30440

   PIN n_30553
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.522 0.163 65.55 ;
      END
   END n_30553

   PIN n_30797
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.114 0.163 56.142 ;
      END
   END n_30797

   PIN n_30876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.026 0.163 63.054 ;
      END
   END n_30876

   PIN n_31014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.002 107.357 14.03 107.52 ;
      END
   END n_31014

   PIN n_31307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.418 0.163 10.446 ;
      END
   END n_31307

   PIN n_31336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.122 107.357 83.15 107.52 ;
      END
   END n_31336

   PIN n_31495
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.482 0.163 10.51 ;
      END
   END n_31495

   PIN n_31518
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.578 107.357 6.606 107.52 ;
      END
   END n_31518

   PIN n_41192
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.106 0.163 37.134 ;
      END
   END n_41192

   PIN n_4674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.45 0.0 30.478 0.163 ;
      END
   END n_4674

   PIN n_4824
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.202 0.0 25.23 0.163 ;
      END
   END n_4824

   PIN n_4835
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.298 0.0 29.326 0.163 ;
      END
   END n_4835

   PIN n_50249
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.234 0.0 21.262 0.163 ;
      END
   END n_50249

   PIN n_50280
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.226 0.163 10.254 ;
      END
   END n_50280

   PIN n_50309
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.666 0.163 7.694 ;
      END
   END n_50309

   PIN n_52277
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.266 0.163 1.294 ;
      END
   END n_52277

   PIN n_55135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 1.202 0.163 1.23 ;
      END
   END n_55135

   PIN n_58287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.522 0.163 1.55 ;
      END
   END n_58287

   PIN n_60578
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.626 0.0 0.654 0.163 ;
      END
   END n_60578

   PIN n_61454
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.53 0.163 44.558 ;
      END
   END n_61454

   PIN n_62185
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.29 0.163 82.318 ;
      END
   END n_62185

   PIN n_62568
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.426 0.163 29.454 ;
      END
   END n_62568

   PIN n_65731
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 17.778 0.163 17.806 ;
      END
   END n_65731

   PIN n_65737
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.714 0.163 17.742 ;
      END
   END n_65737

   PIN n_71280
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.37 0.0 24.398 0.163 ;
      END
   END n_71280

   PIN n_71289
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.354 0.0 18.382 0.163 ;
      END
   END n_71289

   PIN n_95526
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.378 0.0 11.406 0.163 ;
      END
   END n_95526

   PIN n_95541
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.73 0.163 7.758 ;
      END
   END n_95541

   PIN n_97764
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.29 0.163 10.318 ;
      END
   END n_97764

   PIN FE_OFN13766_n_21642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.602 0.0 23.63 0.163 ;
      END
   END FE_OFN13766_n_21642

   PIN FE_OFN17030_n_96760
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.226 0.163 82.254 ;
      END
   END FE_OFN17030_n_96760

   PIN FE_OFN17827_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.93 0.163 90.958 ;
      END
   END FE_OFN17827_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_11_

   PIN FE_OFN17829_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.202 0.163 33.23 ;
      END
   END FE_OFN17829_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_10_

   PIN FE_OFN17831_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.082 0.163 60.11 ;
      END
   END FE_OFN17831_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_9_

   PIN FE_OFN18446_n_30620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.778 0.0 17.806 0.163 ;
      END
   END FE_OFN18446_n_30620

   PIN FE_OFN18448_n_30852
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.242 0.0 16.27 0.163 ;
      END
   END FE_OFN18448_n_30852

   PIN FE_OFN18457_n_27906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.434 0.0 24.462 0.163 ;
      END
   END FE_OFN18457_n_27906

   PIN FE_OFN18870_n_30145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 24.562 99.456 24.59 ;
      END
   END FE_OFN18870_n_30145

   PIN FE_OFN2315_delay_mul_ln34_unr9_unr5_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.346 0.163 79.374 ;
      END
   END FE_OFN2315_delay_mul_ln34_unr9_unr5_stage2_stallmux_z_14_

   PIN FE_OFN2340_delay_mul_ln34_unr9_unr5_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.642 0.163 86.67 ;
      END
   END FE_OFN2340_delay_mul_ln34_unr9_unr5_stage2_stallmux_z_13_

   PIN FE_OFN2342_delay_mul_ln34_unr9_unr5_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 87.986 0.163 88.014 ;
      END
   END FE_OFN2342_delay_mul_ln34_unr9_unr5_stage2_stallmux_z_12_

   PIN FE_OFN271_delay_mul_ln34_unr8_unr5_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.282 0.163 55.31 ;
      END
   END FE_OFN271_delay_mul_ln34_unr8_unr5_stage2_stallmux_z_11_

   PIN FE_OFN273_delay_mul_ln34_unr8_unr5_stage2_stallmux_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.722 0.163 52.75 ;
      END
   END FE_OFN273_delay_mul_ln34_unr8_unr5_stage2_stallmux_z_10_

   PIN FE_OFN275_delay_mul_ln34_unr8_unr5_stage2_stallmux_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.866 0.163 50.894 ;
      END
   END FE_OFN275_delay_mul_ln34_unr8_unr5_stage2_stallmux_z_9_

   PIN FE_OFN287_delay_mul_ln34_unr8_unr5_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.13 0.163 14.158 ;
      END
   END FE_OFN287_delay_mul_ln34_unr8_unr5_stage2_stallmux_z_7_

   PIN FE_OFN6173_n_8289
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 37.106 0.163 37.134 ;
      END
   END FE_OFN6173_n_8289

   PIN FE_OFN6175_n_6867
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.37 0.163 48.398 ;
      END
   END FE_OFN6175_n_6867

   PIN FE_OFN6245_delay_mul_ln34_unr7_unr5_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.674 0.0 2.702 0.163 ;
      END
   END FE_OFN6245_delay_mul_ln34_unr7_unr5_stage2_stallmux_z_14_

   PIN FE_OFN6275_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.274 0.163 52.302 ;
      END
   END FE_OFN6275_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_7_

   PIN FE_OFN6277_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.786 0.163 20.814 ;
      END
   END FE_OFN6277_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_6_

   PIN FE_OFN6279_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.362 0.163 29.39 ;
      END
   END FE_OFN6279_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_5_

   PIN FE_OFN6281_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.618 0.163 21.646 ;
      END
   END FE_OFN6281_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_4_

   PIN FE_OFN6321_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.458 0.163 25.486 ;
      END
   END FE_OFN6321_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_8_

   PIN FE_OFN6326_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 34.546 0.163 34.574 ;
      END
   END FE_OFN6326_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_7_

   PIN FE_OFN6347_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.562 0.163 24.59 ;
      END
   END FE_OFN6347_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_6_

   PIN FE_OFN6350_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.882 0.163 16.91 ;
      END
   END FE_OFN6350_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_5_

   PIN FE_OFN6354_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.298 0.163 29.326 ;
      END
   END FE_OFN6354_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_4_

   PIN FE_OFN6429_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.162 0.163 18.19 ;
      END
   END FE_OFN6429_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_3_

   PIN FE_OFN6431_n_137681
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.882 0.163 40.91 ;
      END
   END FE_OFN6431_n_137681

   PIN FE_OFN6433_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 44.722 0.163 44.75 ;
      END
   END FE_OFN6433_delay_mul_ln34_unr7_unr2_stage2_stallmux_z_2_

   PIN FE_OFN6479_n_137683
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 21.746 0.163 21.774 ;
      END
   END FE_OFN6479_n_137683

   PIN FE_OFN6662_n_41611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.29 0.082 2.318 ;
      END
   END FE_OFN6662_n_41611

   PIN FE_OFN6700_n_41708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.514 0.163 6.542 ;
      END
   END FE_OFN6700_n_41708

   PIN FE_OFN8635_n_31158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.81 0.163 21.838 ;
      END
   END FE_OFN8635_n_31158

   PIN FE_OFN8637_n_31365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.946 0.163 40.974 ;
      END
   END FE_OFN8637_n_31365

   PIN FE_OFN8669_n_30440
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 2.802 99.456 2.83 ;
      END
   END FE_OFN8669_n_30440

   PIN FE_OFN8781_n_22213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.202 0.0 25.23 0.163 ;
      END
   END FE_OFN8781_n_22213

   PIN FE_OFN8824_n_28157
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.626 0.163 40.654 ;
      END
   END FE_OFN8824_n_28157

   PIN FE_OFN8827_n_26678
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.762 0.163 27.79 ;
      END
   END FE_OFN8827_n_26678

   PIN FE_OFN8830_n_26043
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.946 0.163 40.974 ;
      END
   END FE_OFN8830_n_26043

   PIN FE_OFN8832_n_25413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.666 0.163 47.694 ;
      END
   END FE_OFN8832_n_25413

   PIN FE_OFN8942_n_30544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.962 0.163 14.99 ;
      END
   END FE_OFN8942_n_30544

   PIN FE_OFN8993_n_25980
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.002 0.0 30.03 0.163 ;
      END
   END FE_OFN8993_n_25980

   PIN FE_OFN8995_n_26605
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.026 0.0 31.054 0.163 ;
      END
   END FE_OFN8995_n_26605

   PIN FE_OFN8997_n_27189
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.242 0.0 32.27 0.163 ;
      END
   END FE_OFN8997_n_27189

   PIN FE_OFN9000_n_27824
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.394 0.0 33.422 0.163 ;
      END
   END FE_OFN9000_n_27824

   PIN FE_OFN9002_n_28346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.354 0.0 34.382 0.163 ;
      END
   END FE_OFN9002_n_28346

   PIN FE_OFN9004_n_28856
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 35.89 0.0 35.918 0.163 ;
      END
   END FE_OFN9004_n_28856

   PIN FE_OFN9005_n_25363
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.618 0.0 29.646 0.163 ;
      END
   END FE_OFN9005_n_25363

   PIN FE_OFN9008_n_24657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.698 0.0 27.726 0.163 ;
      END
   END FE_OFN9008_n_24657

   PIN FE_OFN9009_n_24023
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 27.698 0.0 27.726 0.163 ;
      END
   END FE_OFN9009_n_24023

   PIN FE_OFN9011_n_23352
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.674 0.0 26.702 0.163 ;
      END
   END FE_OFN9011_n_23352

   PIN FE_OFN9013_n_22755
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.098 0.0 26.126 0.163 ;
      END
   END FE_OFN9013_n_22755

   PIN FE_OFN9015_n_22188
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.306 0.0 24.334 0.163 ;
      END
   END FE_OFN9015_n_22188

   PIN FE_OFN9019_n_21114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.898 0.0 22.926 0.163 ;
      END
   END FE_OFN9019_n_21114

   PIN FE_OFN9021_n_20861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.818 0.0 24.846 0.163 ;
      END
   END FE_OFN9021_n_20861

   PIN FE_OFN9025_n_16099
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.554 0.0 21.582 0.163 ;
      END
   END FE_OFN9025_n_16099

   PIN FE_OFN9031_n_18065
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 83.122 99.456 83.15 ;
      END
   END FE_OFN9031_n_18065

   PIN FE_OFN9051_n_26309
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.674 0.0 18.702 0.163 ;
      END
   END FE_OFN9051_n_26309

   PIN FE_OFN9053_n_26017
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.09 0.0 15.118 0.163 ;
      END
   END FE_OFN9053_n_26017

   PIN FE_OFN9055_n_25387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.258 0.0 14.286 0.163 ;
      END
   END FE_OFN9055_n_25387

   PIN FE_OFN9057_n_24692
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.594 0.0 12.622 0.163 ;
      END
   END FE_OFN9057_n_24692

   PIN FE_OFN9059_n_24066
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.386 0.0 6.414 0.163 ;
      END
   END FE_OFN9059_n_24066

   PIN FE_OFN9061_n_22807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.466 0.0 12.494 0.163 ;
      END
   END FE_OFN9061_n_22807

   PIN FE_OFN9065_n_18510
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.194 0.0 14.222 0.163 ;
      END
   END FE_OFN9065_n_18510

   PIN FE_OFN9227_delay_add_ln34_unr2_unr5_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.002 0.163 30.03 ;
      END
   END FE_OFN9227_delay_add_ln34_unr2_unr5_stage2_stallmux_q_15_

   PIN FE_OFN9455_b_7_9_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 2.162 0.163 2.19 ;
      END
   END FE_OFN9455_b_7_9_1

   PIN FE_OFN9459_b_7_9_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.202 0.163 1.23 ;
      END
   END FE_OFN9459_b_7_9_0

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.09 0.163 79.118 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 88.306 0.163 88.334 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_3_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.346 0.163 71.374 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 61.426 0.163 61.454 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr7_unr2_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 75.506 0.163 75.534 ;
      END
   END delay_mul_ln34_unr7_unr2_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr7_unr2_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.218 0.163 79.246 ;
      END
   END delay_mul_ln34_unr7_unr2_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr7_unr2_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 79.346 0.163 79.374 ;
      END
   END delay_mul_ln34_unr7_unr2_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.626 0.163 48.654 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_10_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 67.826 0.163 67.854 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_11_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.866 0.163 82.894 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.866 0.163 90.894 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.482 0.163 98.51 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.018 0.163 60.046 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.73 0.163 63.758 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_3_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.986 0.163 64.014 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.986 0.163 56.014 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.506 0.163 67.534 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_6_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.442 0.163 67.47 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_7_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 56.946 0.163 56.974 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_8_

   PIN delay_mul_ln34_unr7_unr4_stage2_stallmux_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.186 0.163 75.214 ;
      END
   END delay_mul_ln34_unr7_unr4_stage2_stallmux_z_9_

   PIN delay_mul_ln34_unr7_unr5_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.81 0.0 5.838 0.163 ;
      END
   END delay_mul_ln34_unr7_unr5_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr7_unr5_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.658 0.0 4.686 0.163 ;
      END
   END delay_mul_ln34_unr7_unr5_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.802 0.163 18.83 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.042 0.163 37.07 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.394 0.163 25.422 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr7_unr6_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 29.234 0.163 29.262 ;
      END
   END delay_mul_ln34_unr7_unr6_stage2_stallmux_z_7_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 44.21 99.456 44.238 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 57.842 99.456 57.87 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_11_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 62.962 99.456 62.99 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 34.482 99.456 34.51 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.522 0.163 49.55 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.322 0.163 102.35 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.298 0.163 37.326 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 55.922 99.456 55.95 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_z_10_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 66.162 99.456 66.19 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 71.666 99.456 71.694 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 99.293 45.042 99.456 45.07 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_z_3_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 47.09 99.456 47.118 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 48.242 99.456 48.27 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 54.642 99.456 54.67 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_z_9_

   PIN delay_mul_ln34_unr8_unr2_stage2_stallmux_q_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.562 0.0 40.59 0.163 ;
      END
   END delay_mul_ln34_unr8_unr2_stage2_stallmux_q_10_

   PIN delay_mul_ln34_unr8_unr2_stage2_stallmux_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.466 0.0 44.494 0.163 ;
      END
   END delay_mul_ln34_unr8_unr2_stage2_stallmux_q_11_

   PIN delay_mul_ln34_unr8_unr2_stage2_stallmux_q_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.386 0.0 38.414 0.163 ;
      END
   END delay_mul_ln34_unr8_unr2_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr8_unr2_stage2_stallmux_q_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.274 0.0 36.302 0.163 ;
      END
   END delay_mul_ln34_unr8_unr2_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr8_unr2_stage2_stallmux_q_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.746 0.0 37.774 0.163 ;
      END
   END delay_mul_ln34_unr8_unr2_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr8_unr2_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.514 0.0 30.542 0.163 ;
      END
   END delay_mul_ln34_unr8_unr2_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr8_unr2_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.338 0.0 52.366 0.163 ;
      END
   END delay_mul_ln34_unr8_unr2_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr8_unr2_stage2_stallmux_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.786 0.0 44.814 0.163 ;
      END
   END delay_mul_ln34_unr8_unr2_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr8_unr3_stage2_stallmux_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.562 0.163 40.59 ;
      END
   END delay_mul_ln34_unr8_unr3_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr8_unr3_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 47.602 99.456 47.63 ;
      END
   END delay_mul_ln34_unr8_unr3_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr8_unr3_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 44.722 99.456 44.75 ;
      END
   END delay_mul_ln34_unr8_unr3_stage2_stallmux_z_3_

   PIN delay_mul_ln34_unr8_unr3_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 44.658 99.456 44.686 ;
      END
   END delay_mul_ln34_unr8_unr3_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr8_unr3_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 47.026 99.456 47.054 ;
      END
   END delay_mul_ln34_unr8_unr3_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr8_unr3_stage2_stallmux_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 45.682 99.456 45.71 ;
      END
   END delay_mul_ln34_unr8_unr3_stage2_stallmux_z_6_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.866 0.0 90.894 0.163 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.906 0.163 57.934 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 59.762 99.456 59.79 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 59.122 99.456 59.15 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.65 0.163 25.678 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 17.842 0.163 17.87 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.922 0.163 39.95 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_3_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.842 0.0 17.87 0.163 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.746 107.357 29.774 107.52 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 33.202 99.456 33.23 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr8_unr5_stage2_stallmux_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.242 0.163 48.27 ;
      END
   END delay_mul_ln34_unr8_unr5_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.802 0.0 90.83 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.922 0.0 63.95 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.762 0.0 67.79 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.282 0.0 79.31 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_3_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.218 0.0 79.246 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr8_unr8_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.154 0.0 79.182 0.163 ;
      END
   END delay_mul_ln34_unr8_unr8_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr9_unr5_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.842 0.163 73.87 ;
      END
   END delay_mul_ln34_unr9_unr5_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr9_unr5_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 87.922 0.163 87.95 ;
      END
   END delay_mul_ln34_unr9_unr5_stage2_stallmux_z_11_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.746 0.0 21.774 0.163 ;
      END
   END ispd_clk

   PIN mul_4731_72_n_174
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.41 0.163 71.438 ;
      END
   END mul_4731_72_n_174

   PIN mul_4731_72_n_176
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 83.634 0.163 83.662 ;
      END
   END mul_4731_72_n_176

   PIN n_100254
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.186 0.163 3.214 ;
      END
   END n_100254

   PIN n_104153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 83.762 0.163 83.79 ;
      END
   END n_104153

   PIN n_104383
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 1.138 0.163 1.166 ;
      END
   END n_104383

   PIN n_104960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.45 0.163 6.478 ;
      END
   END n_104960

   PIN n_106245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.138 0.163 1.166 ;
      END
   END n_106245

   PIN n_107448
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.226 0.0 10.254 0.163 ;
      END
   END n_107448

   PIN n_11190
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.978 0.163 37.006 ;
      END
   END n_11190

   PIN n_11199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.282 0.163 71.31 ;
      END
   END n_11199

   PIN n_115952
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.73 0.163 79.758 ;
      END
   END n_115952

   PIN n_116008
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.602 0.163 79.63 ;
      END
   END n_116008

   PIN n_119100
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.698 0.163 67.726 ;
      END
   END n_119100

   PIN n_123852
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.922 0.163 79.95 ;
      END
   END n_123852

   PIN n_137677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 25.586 0.163 25.614 ;
      END
   END n_137677

   PIN n_137679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.914 0.163 36.942 ;
      END
   END n_137679

   PIN n_137732
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 46.962 99.456 46.99 ;
      END
   END n_137732

   PIN n_137734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 43.762 99.456 43.79 ;
      END
   END n_137734

   PIN n_137750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.802 0.163 90.83 ;
      END
   END n_137750

   PIN n_137752
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.722 0.163 20.75 ;
      END
   END n_137752

   PIN n_137754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 30.066 0.163 30.094 ;
      END
   END n_137754

   PIN n_137812
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 40.946 99.456 40.974 ;
      END
   END n_137812

   PIN n_137819
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.21 0.163 52.238 ;
      END
   END n_137819

   PIN n_137834
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.834 0.163 86.862 ;
      END
   END n_137834

   PIN n_137848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.738 0.163 90.766 ;
      END
   END n_137848

   PIN n_137853
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.746 0.163 21.774 ;
      END
   END n_137853

   PIN n_137861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.794 0.163 7.822 ;
      END
   END n_137861

   PIN n_137863
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.754 0.163 40.782 ;
      END
   END n_137863

   PIN n_137869
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 25.522 99.456 25.55 ;
      END
   END n_137869

   PIN n_143924
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.626 0.0 16.654 0.163 ;
      END
   END n_143924

   PIN n_144146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.722 0.163 4.75 ;
      END
   END n_144146

   PIN n_144150
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.066 0.163 6.094 ;
      END
   END n_144150

   PIN n_18035
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.01 0.0 33.038 0.163 ;
      END
   END n_18035

   PIN n_18900
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.226 0.0 2.254 0.163 ;
      END
   END n_18900

   PIN n_19304
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.458 0.0 33.486 0.163 ;
      END
   END n_19304

   PIN n_19335
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.386 0.0 6.414 0.163 ;
      END
   END n_19335

   PIN n_21912
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.098 0.0 34.126 0.163 ;
      END
   END n_21912

   PIN n_22782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.082 0.0 36.11 0.163 ;
      END
   END n_22782

   PIN n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.482 0.163 42.51 ;
      END
   END n_23039

   PIN n_23380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.626 0.0 40.654 0.163 ;
      END
   END n_23380

   PIN n_24049
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.21 0.0 52.238 0.163 ;
      END
   END n_24049

   PIN n_24052
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.482 0.163 34.51 ;
      END
   END n_24052

   PIN n_24067
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.458 0.0 33.486 0.163 ;
      END
   END n_24067

   PIN n_24075
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.514 0.0 6.542 0.163 ;
      END
   END n_24075

   PIN n_24451
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.97 0.0 49.998 0.163 ;
      END
   END n_24451

   PIN n_24681
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.594 0.163 44.622 ;
      END
   END n_24681

   PIN n_24728
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.482 0.0 50.51 0.163 ;
      END
   END n_24728

   PIN n_25378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.034 0.0 2.062 0.163 ;
      END
   END n_25378

   PIN n_25389
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.37 0.0 32.398 0.163 ;
      END
   END n_25389

   PIN n_25428
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.114 0.0 48.142 0.163 ;
      END
   END n_25428

   PIN n_25497
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.498 0.0 80.526 0.163 ;
      END
   END n_25497

   PIN n_26008
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.602 0.163 47.63 ;
      END
   END n_26008

   PIN n_26018
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.474 0.0 31.502 0.163 ;
      END
   END n_26018

   PIN n_26060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.77 0.0 46.798 0.163 ;
      END
   END n_26060

   PIN n_26293
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.202 0.163 49.23 ;
      END
   END n_26293

   PIN n_26654
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.258 0.0 30.286 0.163 ;
      END
   END n_26654

   PIN n_26694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.618 0.0 45.646 0.163 ;
      END
   END n_26694

   PIN n_26911
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.802 0.163 50.83 ;
      END
   END n_26911

   PIN n_27078
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.034 0.0 42.062 0.163 ;
      END
   END n_27078

   PIN n_27222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.802 0.0 90.83 0.163 ;
      END
   END n_27222

   PIN n_27243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 29.554 0.0 29.582 0.163 ;
      END
   END n_27243

   PIN n_27301
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.586 0.163 25.614 ;
      END
   END n_27301

   PIN n_27353
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.058 0.0 43.086 0.163 ;
      END
   END n_27353

   PIN n_27538
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.786 0.163 52.814 ;
      END
   END n_27538

   PIN n_27569
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.85 0.0 28.878 0.163 ;
      END
   END n_27569

   PIN n_27604
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.85 0.0 4.878 0.163 ;
      END
   END n_27604

   PIN n_27697
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.53 0.0 44.558 0.163 ;
      END
   END n_27697

   PIN n_27935
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.178 0.0 40.206 0.163 ;
      END
   END n_27935

   PIN n_28103
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.642 0.163 54.67 ;
      END
   END n_28103

   PIN n_28131
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.266 0.0 25.294 0.163 ;
      END
   END n_28131

   PIN n_28235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.922 0.0 39.95 0.163 ;
      END
   END n_28235

   PIN n_28622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.122 0.163 43.15 ;
      END
   END n_28622

   PIN n_28635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.922 0.163 55.95 ;
      END
   END n_28635

   PIN n_28669
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.394 0.0 25.422 0.163 ;
      END
   END n_28669

   PIN n_29117
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.842 0.163 57.87 ;
      END
   END n_29117

   PIN n_29147
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 21.17 0.0 21.198 0.163 ;
      END
   END n_29147

   PIN n_29434
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.786 0.0 36.814 0.163 ;
      END
   END n_29434

   PIN n_29508
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.53 0.0 12.558 0.163 ;
      END
   END n_29508

   PIN n_29509
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.634 0.0 11.662 0.163 ;
      END
   END n_29509

   PIN n_29548
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.25 0.0 3.278 0.163 ;
      END
   END n_29548

   PIN n_29575
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.37 0.0 8.398 0.163 ;
      END
   END n_29575

   PIN n_29577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.634 0.0 19.662 0.163 ;
      END
   END n_29577

   PIN n_29615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 44.594 99.456 44.622 ;
      END
   END n_29615

   PIN n_29650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.978 0.0 13.006 0.163 ;
      END
   END n_29650

   PIN n_29942
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.242 0.163 64.27 ;
      END
   END n_29942

   PIN n_29972
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.282 0.0 7.31 0.163 ;
      END
   END n_29972

   PIN n_30014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 60.082 99.456 60.11 ;
      END
   END n_30014

   PIN n_30028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 69.362 99.456 69.39 ;
      END
   END n_30028

   PIN n_30271
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.282 0.163 63.31 ;
      END
   END n_30271

   PIN n_30292
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.514 0.0 6.542 0.163 ;
      END
   END n_30292

   PIN n_30345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 82.802 99.456 82.83 ;
      END
   END n_30345

   PIN n_31042
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.293 77.042 99.456 77.07 ;
      END
   END n_31042

   PIN n_31092
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.338 0.0 52.366 0.163 ;
      END
   END n_31092

   PIN n_31487
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.57 0.163 67.598 ;
      END
   END n_31487

   PIN n_42338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.25 0.163 3.278 ;
      END
   END n_42338

   PIN n_42471
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.058 0.163 3.086 ;
      END
   END n_42471

   PIN n_42480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.762 0.163 67.79 ;
      END
   END n_42480

   PIN n_42529
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.082 0.163 68.11 ;
      END
   END n_42529

   PIN n_42530
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.402 0.163 68.43 ;
      END
   END n_42530

   PIN n_42652
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.962 0.163 70.99 ;
      END
   END n_42652

   PIN n_42729
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.266 0.163 73.294 ;
      END
   END n_42729

   PIN n_42730
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.202 0.163 73.23 ;
      END
   END n_42730

   PIN n_42791
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.338 0.163 68.366 ;
      END
   END n_42791

   PIN n_42798
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.234 0.163 37.262 ;
      END
   END n_42798

   PIN n_42801
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 76.082 0.163 76.11 ;
      END
   END n_42801

   PIN n_42843
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.882 0.163 40.91 ;
      END
   END n_42843

   PIN n_42847
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.722 0.163 68.75 ;
      END
   END n_42847

   PIN n_42872
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.17 0.163 37.198 ;
      END
   END n_42872

   PIN n_42953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.026 0.163 79.054 ;
      END
   END n_42953

   PIN n_43001
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 73.33 0.163 73.358 ;
      END
   END n_43001

   PIN n_43074
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.762 0.163 75.79 ;
      END
   END n_43074

   PIN n_43167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.818 0.163 40.846 ;
      END
   END n_43167

   PIN n_43681
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.146 0.163 4.174 ;
      END
   END n_43681

   PIN n_44033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.562 0.163 72.59 ;
      END
   END n_44033

   PIN n_44061
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 72.114 0.163 72.142 ;
      END
   END n_44061

   PIN n_44522
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.922 0.163 71.95 ;
      END
   END n_44522

   PIN n_44523
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 72.37 0.163 72.398 ;
      END
   END n_44523

   PIN n_4772
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.73 0.0 47.758 0.163 ;
      END
   END n_4772

   PIN n_49431
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.778 0.163 17.806 ;
      END
   END n_49431

   PIN n_49913
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.634 0.163 67.662 ;
      END
   END n_49913

   PIN n_50250
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.234 0.0 21.262 0.163 ;
      END
   END n_50250

   PIN n_50281
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.386 0.163 6.414 ;
      END
   END n_50281

   PIN n_50308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 1.074 0.163 1.102 ;
      END
   END n_50308

   PIN n_50379
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.426 0.163 69.454 ;
      END
   END n_50379

   PIN n_50454
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.794 0.163 63.822 ;
      END
   END n_50454

   PIN n_52028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 21.682 0.163 21.71 ;
      END
   END n_52028

   PIN n_52512
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.266 0.163 33.294 ;
      END
   END n_52512

   PIN n_52572
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.082 0.163 4.11 ;
      END
   END n_52572

   PIN n_52708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.01 0.163 41.038 ;
      END
   END n_52708

   PIN n_53209
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.362 0.163 69.39 ;
      END
   END n_53209

   PIN n_54797
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 79.154 0.163 79.182 ;
      END
   END n_54797

   PIN n_54849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.858 0.163 7.886 ;
      END
   END n_54849

   PIN n_54877
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.226 0.163 10.254 ;
      END
   END n_54877

   PIN n_54956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.322 0.163 6.35 ;
      END
   END n_54956

   PIN n_54970
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.098 0.163 10.126 ;
      END
   END n_54970

   PIN n_54980
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.642 0.163 70.67 ;
      END
   END n_54980

   PIN n_55005
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.25 0.163 75.278 ;
      END
   END n_55005

   PIN n_55011
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.106 0.163 77.134 ;
      END
   END n_55011

   PIN n_55098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.034 0.163 10.062 ;
      END
   END n_55098

   PIN n_55101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.45 0.0 22.478 0.163 ;
      END
   END n_55101

   PIN n_55136
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.97 0.0 9.998 0.163 ;
      END
   END n_55136

   PIN n_55151
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.514 0.0 22.542 0.163 ;
      END
   END n_55151

   PIN n_56232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.786 0.163 4.814 ;
      END
   END n_56232

   PIN n_56234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.722 0.163 4.75 ;
      END
   END n_56234

   PIN n_57438
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.034 0.0 18.062 0.163 ;
      END
   END n_57438

   PIN n_57499
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.37 0.0 24.398 0.163 ;
      END
   END n_57499

   PIN n_57501
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.986 0.0 24.014 0.163 ;
      END
   END n_57501

   PIN n_57508
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 6.322 0.0 6.35 0.163 ;
      END
   END n_57508

   PIN n_57682
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 0.946 0.163 0.974 ;
      END
   END n_57682

   PIN n_57709
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 83.57 0.163 83.598 ;
      END
   END n_57709

   PIN n_57710
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 83.506 0.163 83.534 ;
      END
   END n_57710

   PIN n_57792
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.634 0.163 75.662 ;
      END
   END n_57792

   PIN n_57799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 14.002 0.163 14.03 ;
      END
   END n_57799

   PIN n_57875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 9.97 0.163 9.998 ;
      END
   END n_57875

   PIN n_57882
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.002 0.163 6.03 ;
      END
   END n_57882

   PIN n_57917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.034 0.163 10.062 ;
      END
   END n_57917

   PIN n_58050
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.898 0.163 70.926 ;
      END
   END n_58050

   PIN n_58096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 1.586 0.163 1.614 ;
      END
   END n_58096

   PIN n_58458
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.162 0.163 10.19 ;
      END
   END n_58458

   PIN n_58653
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 0.882 0.163 0.91 ;
      END
   END n_58653

   PIN n_58825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.162 0.163 74.19 ;
      END
   END n_58825

   PIN n_58842
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 52.402 0.163 52.43 ;
      END
   END n_58842

   PIN n_58893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 83.698 0.163 83.726 ;
      END
   END n_58893

   PIN n_58929
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.442 0.163 3.47 ;
      END
   END n_58929

   PIN n_58997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.354 0.0 10.382 0.163 ;
      END
   END n_58997

   PIN n_58998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.714 0.0 17.742 0.163 ;
      END
   END n_58998

   PIN n_59262
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.162 0.163 10.19 ;
      END
   END n_59262

   PIN n_59928
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.186 0.0 19.214 0.163 ;
      END
   END n_59928

   PIN n_60313
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.85 0.0 20.878 0.163 ;
      END
   END n_60313

   PIN n_60331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.738 0.0 18.766 0.163 ;
      END
   END n_60331

   PIN n_60641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.706 0.163 6.734 ;
      END
   END n_60641

   PIN n_60716
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 83.442 0.163 83.47 ;
      END
   END n_60716

   PIN n_60751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 6.642 0.163 6.67 ;
      END
   END n_60751

   PIN n_61044
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 0.946 0.163 0.974 ;
      END
   END n_61044

   PIN n_61084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.906 0.0 9.934 0.163 ;
      END
   END n_61084

   PIN n_61701
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.098 0.163 10.126 ;
      END
   END n_61701

   PIN n_62186
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.162 0.163 82.19 ;
      END
   END n_62186

   PIN n_62600
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.354 0.163 10.382 ;
      END
   END n_62600

   PIN n_62607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.29 0.163 10.318 ;
      END
   END n_62607

   PIN n_63108
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.522 0.0 1.55 0.163 ;
      END
   END n_63108

   PIN n_63353
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.45 0.0 14.478 0.163 ;
      END
   END n_63353

   PIN n_63538
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.938 0.163 77.966 ;
      END
   END n_63538

   PIN n_63691
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.69 0.163 40.718 ;
      END
   END n_63691

   PIN n_65307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.874 0.163 13.902 ;
      END
   END n_65307

   PIN n_6646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.49 0.0 29.518 0.163 ;
      END
   END n_6646

   PIN n_71288
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.418 0.0 18.446 0.163 ;
      END
   END n_71288

   PIN n_71418
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.066 0.163 14.094 ;
      END
   END n_71418

   PIN n_71433
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 14.002 0.163 14.03 ;
      END
   END n_71433

   PIN n_7178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.138 0.163 33.166 ;
      END
   END n_7178

   PIN n_71966
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.554 0.163 21.582 ;
      END
   END n_71966

   PIN n_81058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.314 0.0 19.342 0.163 ;
      END
   END n_81058

   PIN n_8266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.242 0.163 16.27 ;
      END
   END n_8266

   PIN n_83289
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.642 0.0 14.67 0.163 ;
      END
   END n_83289

   PIN n_83679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.562 0.0 16.59 0.163 ;
      END
   END n_83679

   PIN n_8374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.242 0.163 32.27 ;
      END
   END n_8374

   PIN n_8393
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.85 0.163 36.878 ;
      END
   END n_8393

   PIN n_85475
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.426 0.0 13.454 0.163 ;
      END
   END n_85475

   PIN n_85700
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.922 0.163 7.95 ;
      END
   END n_85700

   PIN n_85705
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 7.922 0.163 7.95 ;
      END
   END n_85705

   PIN n_89145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.474 0.0 15.502 0.163 ;
      END
   END n_89145

   PIN n_89166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.45 0.0 14.478 0.163 ;
      END
   END n_89166

   PIN n_89167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.706 0.0 14.734 0.163 ;
      END
   END n_89167

   PIN n_91981
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.602 0.163 7.63 ;
      END
   END n_91981

   PIN n_92794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 1.01 0.163 1.038 ;
      END
   END n_92794

   PIN n_92795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.738 0.0 10.766 0.163 ;
      END
   END n_92795

   PIN n_94774
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.754 0.0 0.782 0.163 ;
      END
   END n_94774

   PIN n_94777
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.69 0.0 0.718 0.163 ;
      END
   END n_94777

   PIN n_95516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.49 0.0 13.518 0.163 ;
      END
   END n_95516

   PIN n_95527
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.762 0.0 11.79 0.163 ;
      END
   END n_95527

   PIN n_95530
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.826 0.0 11.854 0.163 ;
      END
   END n_95530

   PIN n_95531
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 6.45 0.0 6.478 0.163 ;
      END
   END n_95531

   PIN n_95538
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.074 0.163 1.102 ;
      END
   END n_95538

   PIN n_95542
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 1.01 0.163 1.038 ;
      END
   END n_95542

   PIN n_97281
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.778 0.0 25.806 0.163 ;
      END
   END n_97281

   PIN n_97761
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 13.938 0.163 13.966 ;
      END
   END n_97761

   PIN n_99215
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.698 0.0 11.726 0.163 ;
      END
   END n_99215

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 99.456 107.52 ;
      LAYER V1 ;
         RECT 0.0 0.0 99.456 107.52 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 99.456 107.52 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 99.456 107.52 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 99.456 107.52 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 99.456 107.52 ;
      LAYER M1 ;
         RECT 0.0 0.0 99.456 107.52 ;
   END
END h8_mgc_matrix_mult_b

MACRO h7_mgc_matrix_mult_b
   CLASS BLOCK ;
   FOREIGN h7 ;
   ORIGIN 0 0 ;
   SIZE 137.792 BY 36.48 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN15487_FE_OFN12404_n_112269
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.498 36.317 104.526 36.48 ;
      END
   END FE_OCPN15487_FE_OFN12404_n_112269

   PIN FE_OCPN15496_FE_OFN13305_n_143019
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.242 36.317 112.27 36.48 ;
      END
   END FE_OCPN15496_FE_OFN13305_n_143019

   PIN FE_OCPN15502_n_111893
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.53 36.317 108.558 36.48 ;
      END
   END FE_OCPN15502_n_111893

   PIN FE_OCPN15568_FE_OFN11385_n_210
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.666 36.317 119.694 36.48 ;
      END
   END FE_OCPN15568_FE_OFN11385_n_210

   PIN FE_OCPN15572_FE_OFN12407_n_143087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.146 36.317 100.174 36.48 ;
      END
   END FE_OCPN15572_FE_OFN12407_n_143087

   PIN FE_OCPN15750_FE_OFN13746_n_143074
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.914 36.317 108.942 36.48 ;
      END
   END FE_OCPN15750_FE_OFN13746_n_143074

   PIN FE_OFN10392_b_1_1_6
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.866 36.317 114.894 36.48 ;
      END
   END FE_OFN10392_b_1_1_6

   PIN FE_OFN10397_b_1_1_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.082 36.317 116.11 36.48 ;
      END
   END FE_OFN10397_b_1_1_4

   PIN FE_OFN10398_b_1_1_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.154 36.317 119.182 36.48 ;
      END
   END FE_OFN10398_b_1_1_4

   PIN FE_OFN10400_b_1_1_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.01 36.317 113.038 36.48 ;
      END
   END FE_OFN10400_b_1_1_3

   PIN FE_OFN10402_b_1_1_2
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 118.258 36.398 118.286 36.48 ;
      END
   END FE_OFN10402_b_1_1_2

   PIN FE_OFN10409_b_1_1_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.162 36.398 106.19 36.48 ;
      END
   END FE_OFN10409_b_1_1_0

   PIN FE_OFN11381_n_142891
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.922 36.317 103.95 36.48 ;
      END
   END FE_OFN11381_n_142891

   PIN FE_OFN11476_n_143637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.674 36.317 130.702 36.48 ;
      END
   END FE_OFN11476_n_143637

   PIN FE_OFN11985_n_143017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.634 36.317 123.662 36.48 ;
      END
   END FE_OFN11985_n_143017

   PIN FE_OFN11987_n_143017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.666 36.317 127.694 36.48 ;
      END
   END FE_OFN11987_n_143017

   PIN FE_OFN11988_n_143017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 33.714 137.792 33.742 ;
      END
   END FE_OFN11988_n_143017

   PIN FE_OFN12353_n_112222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.01 36.317 105.038 36.48 ;
      END
   END FE_OFN12353_n_112222

   PIN FE_OFN12404_n_112269
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.41 36.317 111.438 36.48 ;
      END
   END FE_OFN12404_n_112269

   PIN FE_OFN12662_n_142936
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.218 36.317 119.246 36.48 ;
      END
   END FE_OFN12662_n_142936

   PIN FE_OFN12694_n_142879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.17 36.317 109.198 36.48 ;
      END
   END FE_OFN12694_n_142879

   PIN FE_OFN12697_n_142879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.85 36.317 108.878 36.48 ;
      END
   END FE_OFN12697_n_142879

   PIN FE_OFN12701_n_142878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.426 36.317 109.454 36.48 ;
      END
   END FE_OFN12701_n_142878

   PIN FE_OFN12702_n_142878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.298 36.317 109.326 36.48 ;
      END
   END FE_OFN12702_n_142878

   PIN FE_OFN12703_n_142878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.346 36.317 111.374 36.48 ;
      END
   END FE_OFN12703_n_142878

   PIN FE_OFN12708_n_142877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.954 36.317 107.982 36.48 ;
      END
   END FE_OFN12708_n_142877

   PIN FE_OFN12741_n_143073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.442 36.317 131.47 36.48 ;
      END
   END FE_OFN12741_n_143073

   PIN FE_OFN12742_n_143073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.266 36.317 89.294 36.48 ;
      END
   END FE_OFN12742_n_143073

   PIN FE_OFN13304_n_143019
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.106 36.317 117.134 36.48 ;
      END
   END FE_OFN13304_n_143019

   PIN FE_OFN13307_n_143018
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.45 36.317 118.478 36.48 ;
      END
   END FE_OFN13307_n_143018

   PIN FE_OFN13496_n_111726
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 124.978 36.317 125.006 36.48 ;
      END
   END FE_OFN13496_n_111726

   PIN FE_OFN13571_n_143090
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.37 36.317 104.398 36.48 ;
      END
   END FE_OFN13571_n_143090

   PIN FE_OFN13575_n_143090
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.434 36.317 96.462 36.48 ;
      END
   END FE_OFN13575_n_143090

   PIN FE_OFN13593_n_142824
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.794 36.317 111.822 36.48 ;
      END
   END FE_OFN13593_n_142824

   PIN FE_OFN13605_n_142822
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.274 36.317 116.302 36.48 ;
      END
   END FE_OFN13605_n_142822

   PIN FE_OFN13648_n_143638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.258 36.317 118.286 36.48 ;
      END
   END FE_OFN13648_n_143638

   PIN FE_OFN13649_n_143638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.218 36.317 119.246 36.48 ;
      END
   END FE_OFN13649_n_143638

   PIN FE_OFN14250_n_140259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.506 36.317 131.534 36.48 ;
      END
   END FE_OFN14250_n_140259

   PIN FE_OFN14252_n_140259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.962 36.317 118.99 36.48 ;
      END
   END FE_OFN14252_n_140259

   PIN FE_OFN14255_n_140259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.642 36.317 118.67 36.48 ;
      END
   END FE_OFN14255_n_140259

   PIN FE_OFN14256_n_140259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.658 36.317 116.686 36.48 ;
      END
   END FE_OFN14256_n_140259

   PIN FE_OFN14257_n_140259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.538 36.317 127.566 36.48 ;
      END
   END FE_OFN14257_n_140259

   PIN FE_OFN14259_n_140259
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.466 36.317 116.494 36.48 ;
      END
   END FE_OFN14259_n_140259

   PIN FE_OFN14394_n_142835
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.122 36.317 115.15 36.48 ;
      END
   END FE_OFN14394_n_142835

   PIN FE_OFN14886_n_590
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.41 36.317 119.438 36.48 ;
      END
   END FE_OFN14886_n_590

   PIN FE_OFN15897_n_143087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.266 36.317 121.294 36.48 ;
      END
   END FE_OFN15897_n_143087

   PIN FE_OFN16418_b_1_1_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.002 36.317 110.03 36.48 ;
      END
   END FE_OFN16418_b_1_1_3

   PIN FE_OFN16622_delay_add_ln34_unr2_unr9_stage2_stallmux_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.866 36.317 2.894 36.48 ;
      END
   END FE_OFN16622_delay_add_ln34_unr2_unr9_stage2_stallmux_z_14_

   PIN FE_OFN16914_n_19194
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.642 0.0 54.67 0.163 ;
      END
   END FE_OFN16914_n_19194

   PIN FE_OFN17087_n_142823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.442 36.317 123.47 36.48 ;
      END
   END FE_OFN17087_n_142823

   PIN FE_OFN17137_n_15473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 131.506 36.317 131.534 36.48 ;
      END
   END FE_OFN17137_n_15473

   PIN FE_OFN18629_b_1_1_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.106 36.317 109.134 36.48 ;
      END
   END FE_OFN18629_b_1_1_5

   PIN FE_OFN18763_n_142881
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.29 36.317 106.318 36.48 ;
      END
   END FE_OFN18763_n_142881

   PIN FE_OFN18849_n_142838
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.93 36.317 114.958 36.48 ;
      END
   END FE_OFN18849_n_142838

   PIN FE_OFN1973_n_17469
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.698 36.317 123.726 36.48 ;
      END
   END FE_OFN1973_n_17469

   PIN FE_OFN2297_n_142894
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.994 36.317 115.022 36.48 ;
      END
   END FE_OFN2297_n_142894

   PIN FE_OFN2689_n_142837
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.21 36.317 100.238 36.48 ;
      END
   END FE_OFN2689_n_142837

   PIN FE_OFN2744_n_123691
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.498 36.317 96.526 36.48 ;
      END
   END FE_OFN2744_n_123691

   PIN FE_OFN2832_n_142934
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.73 36.317 119.758 36.48 ;
      END
   END FE_OFN2832_n_142934

   PIN FE_OFN2833_n_142934
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.602 36.317 127.63 36.48 ;
      END
   END FE_OFN2833_n_142934

   PIN FE_OFN2851_n_111724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.282 36.317 135.31 36.48 ;
      END
   END FE_OFN2851_n_111724

   PIN delay_add_ln34_unr2_unr4_stage2_stallmux_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.89 36.317 11.918 36.48 ;
      END
   END delay_add_ln34_unr2_unr4_stage2_stallmux_q_0_

   PIN delay_add_ln34_unr2_unr4_stage2_stallmux_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.266 36.317 17.294 36.48 ;
      END
   END delay_add_ln34_unr2_unr4_stage2_stallmux_q_1_

   PIN delay_add_ln34_unr2_unr4_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.378 36.317 19.406 36.48 ;
      END
   END delay_add_ln34_unr2_unr4_stage2_stallmux_q_2_

   PIN delay_add_ln34_unr2_unr4_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.866 36.317 18.894 36.48 ;
      END
   END delay_add_ln34_unr2_unr4_stage2_stallmux_q_3_

   PIN delay_add_ln34_unr2_unr4_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.562 36.317 8.59 36.48 ;
      END
   END delay_add_ln34_unr2_unr4_stage2_stallmux_q_4_

   PIN delay_add_ln34_unr2_unr4_stage2_stallmux_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.578 36.317 14.606 36.48 ;
      END
   END delay_add_ln34_unr2_unr4_stage2_stallmux_q_5_

   PIN delay_add_ln34_unr2_unr4_stage2_stallmux_q_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.562 36.317 8.59 36.48 ;
      END
   END delay_add_ln34_unr2_unr4_stage2_stallmux_q_6_

   PIN delay_add_ln34_unr2_unr4_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.186 36.317 3.214 36.48 ;
      END
   END delay_add_ln34_unr2_unr4_stage2_stallmux_q_7_

   PIN mul_4376_72_n_153
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.066 36.317 102.094 36.48 ;
      END
   END mul_4376_72_n_153

   PIN mul_4376_72_n_154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.074 36.317 105.102 36.48 ;
      END
   END mul_4376_72_n_154

   PIN mul_4376_72_n_275
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.658 36.317 116.686 36.48 ;
      END
   END mul_4376_72_n_275

   PIN mul_4376_72_n_282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.17 36.317 117.198 36.48 ;
      END
   END mul_4376_72_n_282

   PIN mul_4376_72_n_287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.674 36.317 122.702 36.48 ;
      END
   END mul_4376_72_n_287

   PIN mul_4376_72_n_288
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.33 36.317 121.358 36.48 ;
      END
   END mul_4376_72_n_288

   PIN mul_4376_72_n_290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.442 36.317 115.47 36.48 ;
      END
   END mul_4376_72_n_290

   PIN mul_4379_72_n_336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.178 36.317 104.206 36.48 ;
      END
   END mul_4379_72_n_336

   PIN mul_4384_72_n_309
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.69 36.317 120.718 36.48 ;
      END
   END mul_4384_72_n_309

   PIN mul_4385_72_n_188
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.754 36.317 104.782 36.48 ;
      END
   END mul_4385_72_n_188

   PIN mul_4385_72_n_196
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.834 36.317 102.862 36.48 ;
      END
   END mul_4385_72_n_196

   PIN mul_4385_72_n_197
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.354 36.317 98.382 36.48 ;
      END
   END mul_4385_72_n_197

   PIN mul_4385_72_n_198
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.986 36.317 104.014 36.48 ;
      END
   END mul_4385_72_n_198

   PIN mul_4385_72_n_226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.418 36.317 106.446 36.48 ;
      END
   END mul_4385_72_n_226

   PIN mul_4385_72_n_228
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.562 36.317 96.59 36.48 ;
      END
   END mul_4385_72_n_228

   PIN mul_4385_72_n_253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.594 36.317 92.622 36.48 ;
      END
   END mul_4385_72_n_253

   PIN mul_4385_72_n_258
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.674 36.317 98.702 36.48 ;
      END
   END mul_4385_72_n_258

   PIN mul_4385_72_n_291
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.826 36.317 115.854 36.48 ;
      END
   END mul_4385_72_n_291

   PIN mul_4385_72_n_293
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.202 36.317 89.23 36.48 ;
      END
   END mul_4385_72_n_293

   PIN mul_4385_72_n_297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.786 36.317 92.814 36.48 ;
      END
   END mul_4385_72_n_297

   PIN n_111895
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.25 36.317 115.278 36.48 ;
      END
   END n_111895

   PIN n_112002
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.914 36.317 116.942 36.48 ;
      END
   END n_112002

   PIN n_112222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.194 36.398 102.222 36.48 ;
      END
   END n_112222

   PIN n_114682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.874 36.317 109.902 36.48 ;
      END
   END n_114682

   PIN n_114776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.282 36.317 111.31 36.48 ;
      END
   END n_114776

   PIN n_114795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.242 36.317 120.27 36.48 ;
      END
   END n_114795

   PIN n_115233
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.714 36.317 121.742 36.48 ;
      END
   END n_115233

   PIN n_115252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.434 36.317 96.462 36.48 ;
      END
   END n_115252

   PIN n_115271
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.754 36.317 120.782 36.48 ;
      END
   END n_115271

   PIN n_115828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.738 36.317 90.766 36.48 ;
      END
   END n_115828

   PIN n_116358
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.33 36.317 113.358 36.48 ;
      END
   END n_116358

   PIN n_116509
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.202 36.317 113.23 36.48 ;
      END
   END n_116509

   PIN n_116701
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.818 36.317 112.846 36.48 ;
      END
   END n_116701

   PIN n_116804
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.266 36.317 113.294 36.48 ;
      END
   END n_116804

   PIN n_116835
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.074 36.317 113.102 36.48 ;
      END
   END n_116835

   PIN n_118255
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.474 36.317 95.502 36.48 ;
      END
   END n_118255

   PIN n_118393
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.834 36.317 102.862 36.48 ;
      END
   END n_118393

   PIN n_118706
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.434 36.317 112.462 36.48 ;
      END
   END n_118706

   PIN n_120518
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.498 36.317 112.526 36.48 ;
      END
   END n_120518

   PIN n_121402
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.882 36.317 104.91 36.48 ;
      END
   END n_121402

   PIN n_121961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.386 36.317 94.414 36.48 ;
      END
   END n_121961

   PIN n_122290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.17 36.317 109.198 36.48 ;
      END
   END n_122290

   PIN n_122291
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.298 36.317 109.326 36.48 ;
      END
   END n_122291

   PIN n_122325
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.234 36.317 109.262 36.48 ;
      END
   END n_122325

   PIN n_122457
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.794 36.317 103.822 36.48 ;
      END
   END n_122457

   PIN n_123073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.002 36.317 94.03 36.48 ;
      END
   END n_123073

   PIN n_123201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.138 36.317 113.166 36.48 ;
      END
   END n_123201

   PIN n_123230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.882 36.317 112.91 36.48 ;
      END
   END n_123230

   PIN n_123532
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.69 36.317 96.718 36.48 ;
      END
   END n_123532

   PIN n_123533
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.306 36.317 96.334 36.48 ;
      END
   END n_123533

   PIN n_123541
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.69 36.317 96.718 36.48 ;
      END
   END n_123541

   PIN n_123699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.258 36.317 94.286 36.48 ;
      END
   END n_123699

   PIN n_123707
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.826 36.317 99.854 36.48 ;
      END
   END n_123707

   PIN n_123732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.986 36.317 96.014 36.48 ;
      END
   END n_123732

   PIN n_124236
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.786 36.317 108.814 36.48 ;
      END
   END n_124236

   PIN n_124424
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.01 36.317 89.038 36.48 ;
      END
   END n_124424

   PIN n_124618
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.562 36.317 96.59 36.48 ;
      END
   END n_124618

   PIN n_124619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.114 36.317 96.142 36.48 ;
      END
   END n_124619

   PIN n_124704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.066 36.317 94.094 36.48 ;
      END
   END n_124704

   PIN n_124724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.13 36.317 94.158 36.48 ;
      END
   END n_124724

   PIN n_124900
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.058 36.317 99.086 36.48 ;
      END
   END n_124900

   PIN n_124901
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.378 36.317 99.406 36.48 ;
      END
   END n_124901

   PIN n_125656
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.538 36.317 103.566 36.48 ;
      END
   END n_125656

   PIN n_125817
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.322 36.317 94.35 36.48 ;
      END
   END n_125817

   PIN n_127134
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.602 36.317 95.63 36.48 ;
      END
   END n_127134

   PIN n_127158
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.682 36.317 101.71 36.48 ;
      END
   END n_127158

   PIN n_127272
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.85 36.317 92.878 36.48 ;
      END
   END n_127272

   PIN n_127322
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.082 36.317 100.11 36.48 ;
      END
   END n_127322

   PIN n_127852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.914 36.317 92.942 36.48 ;
      END
   END n_127852

   PIN n_127963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.074 36.317 89.102 36.48 ;
      END
   END n_127963

   PIN n_128562
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.754 36.317 96.782 36.48 ;
      END
   END n_128562

   PIN n_128563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.978 36.317 93.006 36.48 ;
      END
   END n_128563

   PIN n_128827
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.802 36.317 98.83 36.48 ;
      END
   END n_128827

   PIN n_128963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.138 36.317 89.166 36.48 ;
      END
   END n_128963

   PIN n_129001
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.202 36.317 89.23 36.48 ;
      END
   END n_129001

   PIN n_129914
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.114 36.317 104.142 36.48 ;
      END
   END n_129914

   PIN n_131586
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.362 36.317 85.39 36.48 ;
      END
   END n_131586

   PIN n_131938
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.538 36.317 119.566 36.48 ;
      END
   END n_131938

   PIN n_142879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.354 36.317 106.382 36.48 ;
      END
   END n_142879

   PIN n_142933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.322 36.317 102.35 36.48 ;
      END
   END n_142933

   PIN n_142934
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.882 36.398 96.91 36.48 ;
      END
   END n_142934

   PIN n_142935
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.522 36.317 113.55 36.48 ;
      END
   END n_142935

   PIN n_143076
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.594 36.317 108.622 36.48 ;
      END
   END n_143076

   PIN n_143077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.578 36.317 102.606 36.48 ;
      END
   END n_143077

   PIN n_143794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.042 36.317 93.07 36.48 ;
      END
   END n_143794

   PIN n_143845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.642 36.317 102.67 36.48 ;
      END
   END n_143845

   PIN n_16174
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 5.042 137.792 5.07 ;
      END
   END n_16174

   PIN n_16223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.426 36.317 109.454 36.48 ;
      END
   END n_16223

   PIN n_16370
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.938 36.317 109.966 36.48 ;
      END
   END n_16370

   PIN n_16624
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.218 36.317 111.246 36.48 ;
      END
   END n_16624

   PIN n_17775
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.362 36.317 109.39 36.48 ;
      END
   END n_17775

   PIN n_18083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.474 36.317 111.502 36.48 ;
      END
   END n_18083

   PIN n_19629
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.082 0.0 20.11 0.163 ;
      END
   END n_19629

   PIN n_2592
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.97 36.317 121.998 36.48 ;
      END
   END n_2592

   PIN n_31935
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.018 36.317 116.046 36.48 ;
      END
   END n_31935

   PIN n_32008
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.73 36.317 111.758 36.48 ;
      END
   END n_32008

   PIN n_32014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.786 36.317 108.814 36.48 ;
      END
   END n_32014

   PIN n_32066
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.642 36.317 110.67 36.48 ;
      END
   END n_32066

   PIN n_32240
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.602 36.317 111.63 36.48 ;
      END
   END n_32240

   PIN n_32283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.21 36.317 116.238 36.48 ;
      END
   END n_32283

   PIN n_32342
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.474 36.317 111.502 36.48 ;
      END
   END n_32342

   PIN n_32407
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.082 36.317 108.11 36.48 ;
      END
   END n_32407

   PIN n_32494
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.05 36.317 104.078 36.48 ;
      END
   END n_32494

   PIN n_32869
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.106 36.317 93.134 36.48 ;
      END
   END n_32869

   PIN n_32877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.722 36.317 92.75 36.48 ;
      END
   END n_32877

   PIN n_33394
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.722 36.317 116.75 36.48 ;
      END
   END n_33394

   PIN n_33847
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.994 36.317 107.022 36.48 ;
      END
   END n_33847

   PIN n_34034
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.89 36.317 99.918 36.48 ;
      END
   END n_34034

   PIN n_34107
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.978 36.317 109.006 36.48 ;
      END
   END n_34107

   PIN n_34672
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.666 36.317 111.694 36.48 ;
      END
   END n_34672

   PIN n_34854
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.042 36.317 109.07 36.48 ;
      END
   END n_34854

   PIN n_34945
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.138 36.317 105.166 36.48 ;
      END
   END n_34945

   PIN n_35146
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.538 36.317 111.566 36.48 ;
      END
   END n_35146

   PIN n_35659
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.242 36.317 104.27 36.48 ;
      END
   END n_35659

   PIN n_35677
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.578 36.317 94.606 36.48 ;
      END
   END n_35677

   PIN n_35915
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.002 36.317 102.03 36.48 ;
      END
   END n_35915

   PIN n_35916
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.402 36.317 100.43 36.48 ;
      END
   END n_35916

   PIN n_36035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.642 36.317 94.67 36.48 ;
      END
   END n_36035

   PIN n_36226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.65 36.317 97.678 36.48 ;
      END
   END n_36226

   PIN n_36445
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.554 36.317 93.582 36.48 ;
      END
   END n_36445

   PIN n_36448
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.162 36.317 98.19 36.48 ;
      END
   END n_36448

   PIN n_36459
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.85 36.317 92.878 36.48 ;
      END
   END n_36459

   PIN n_36620
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.17 36.317 93.198 36.48 ;
      END
   END n_36620

   PIN n_36625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.658 36.317 92.686 36.48 ;
      END
   END n_36625

   PIN n_36656
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.394 36.317 97.422 36.48 ;
      END
   END n_36656

   PIN n_47622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.466 36.317 100.494 36.48 ;
      END
   END n_47622

   PIN n_47691
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.146 36.317 100.174 36.48 ;
      END
   END n_47691

   PIN n_48142
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.906 36.317 97.934 36.48 ;
      END
   END n_48142

   PIN n_49325
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.626 36.317 96.654 36.48 ;
      END
   END n_49325

   PIN n_49408
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.482 36.317 98.51 36.48 ;
      END
   END n_49408

   PIN n_49409
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.546 36.317 98.574 36.48 ;
      END
   END n_49409

   PIN n_4967
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.706 36.317 110.734 36.48 ;
      END
   END n_4967

   PIN n_58898
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.81 36.317 117.838 36.48 ;
      END
   END n_58898

   PIN n_64452
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.978 36.317 117.006 36.48 ;
      END
   END n_64452

   PIN n_64453
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.146 36.317 116.174 36.48 ;
      END
   END n_64453

   PIN n_7726
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 24.306 137.792 24.334 ;
      END
   END n_7726

   PIN FE_OCPN15495_n_143017
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.762 36.317 123.79 36.48 ;
      END
   END FE_OCPN15495_n_143017

   PIN FE_OCPN15497_FE_OFN13305_n_143019
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.794 36.317 111.822 36.48 ;
      END
   END FE_OCPN15497_FE_OFN13305_n_143019

   PIN FE_OCPN15516_FE_OFN13305_n_143019
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.986 36.317 104.014 36.48 ;
      END
   END FE_OCPN15516_FE_OFN13305_n_143019

   PIN FE_OCPN15545_n_143577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.058 36.317 115.086 36.48 ;
      END
   END FE_OCPN15545_n_143577

   PIN FE_OCPN15594_FE_OFN11474_n_143637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.954 36.317 115.982 36.48 ;
      END
   END FE_OCPN15594_FE_OFN11474_n_143637

   PIN FE_OCPN15605_n_142891
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.85 36.317 116.878 36.48 ;
      END
   END FE_OCPN15605_n_142891

   PIN FE_OCPN15647_n_142835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.41 36.317 119.438 36.48 ;
      END
   END FE_OCPN15647_n_142835

   PIN FE_OCPN15669_FE_OFN13856_n_142821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.618 36.317 101.646 36.48 ;
      END
   END FE_OCPN15669_FE_OFN13856_n_142821

   PIN FE_OFN10378_b_1_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.13 36.317 102.158 36.48 ;
      END
   END FE_OFN10378_b_1_4_1

   PIN FE_OFN10380_b_1_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.378 36.317 115.406 36.48 ;
      END
   END FE_OFN10380_b_1_4_0

   PIN FE_OFN10407_b_1_1_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.53 36.317 116.558 36.48 ;
      END
   END FE_OFN10407_b_1_1_1

   PIN FE_OFN10408_b_1_1_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.458 36.317 105.486 36.48 ;
      END
   END FE_OFN10408_b_1_1_0

   PIN FE_OFN10414_b_1_0_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.834 36.317 110.862 36.48 ;
      END
   END FE_OFN10414_b_1_0_7

   PIN FE_OFN10416_b_1_0_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.698 36.317 99.726 36.48 ;
      END
   END FE_OFN10416_b_1_0_5

   PIN FE_OFN10420_b_1_0_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.266 36.317 105.294 36.48 ;
      END
   END FE_OFN10420_b_1_0_3

   PIN FE_OFN10424_b_1_0_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.97 36.317 97.998 36.48 ;
      END
   END FE_OFN10424_b_1_0_0

   PIN FE_OFN11379_n_142891
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.858 36.317 103.886 36.48 ;
      END
   END FE_OFN11379_n_142891

   PIN FE_OFN11389_n_210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.522 36.317 121.55 36.48 ;
      END
   END FE_OFN11389_n_210

   PIN FE_OFN11473_n_143637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.738 36.317 130.766 36.48 ;
      END
   END FE_OFN11473_n_143637

   PIN FE_OFN11539_n_111724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.978 36.317 117.006 36.48 ;
      END
   END FE_OFN11539_n_111724

   PIN FE_OFN11540_n_111724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.602 36.317 119.63 36.48 ;
      END
   END FE_OFN11540_n_111724

   PIN FE_OFN11952_n_143577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.09 36.317 119.118 36.48 ;
      END
   END FE_OFN11952_n_143577

   PIN FE_OFN11983_n_143017
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.514 36.317 118.542 36.48 ;
      END
   END FE_OFN11983_n_143017

   PIN FE_OFN12403_n_112269
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 127.666 36.317 127.694 36.48 ;
      END
   END FE_OFN12403_n_112269

   PIN FE_OFN12406_n_143087
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.042 36.317 117.07 36.48 ;
      END
   END FE_OFN12406_n_143087

   PIN FE_OFN12407_n_143087
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.77 36.317 110.798 36.48 ;
      END
   END FE_OFN12407_n_143087

   PIN FE_OFN12658_n_142936
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.698 36.317 115.726 36.48 ;
      END
   END FE_OFN12658_n_142936

   PIN FE_OFN12659_n_142936
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.77 36.317 110.798 36.48 ;
      END
   END FE_OFN12659_n_142936

   PIN FE_OFN12669_n_142934
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.874 36.317 117.902 36.48 ;
      END
   END FE_OFN12669_n_142934

   PIN FE_OFN12678_n_142893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.442 36.317 107.47 36.48 ;
      END
   END FE_OFN12678_n_142893

   PIN FE_OFN12691_n_142880
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 124.21 36.317 124.238 36.48 ;
      END
   END FE_OFN12691_n_142880

   PIN FE_OFN12705_n_142877
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.914 36.317 108.942 36.48 ;
      END
   END FE_OFN12705_n_142877

   PIN FE_OFN12740_n_143073
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 33.778 137.792 33.806 ;
      END
   END FE_OFN12740_n_143073

   PIN FE_OFN12748_n_143115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.85 36.398 116.878 36.48 ;
      END
   END FE_OFN12748_n_143115

   PIN FE_OFN13299_n_143020
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.674 36.317 106.702 36.48 ;
      END
   END FE_OFN13299_n_143020

   PIN FE_OFN13305_n_143019
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.37 36.317 112.398 36.48 ;
      END
   END FE_OFN13305_n_143019

   PIN FE_OFN13311_n_143018
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 122.034 36.317 122.062 36.48 ;
      END
   END FE_OFN13311_n_143018

   PIN FE_OFN13320_n_142976
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.474 36.317 119.502 36.48 ;
      END
   END FE_OFN13320_n_142976

   PIN FE_OFN13322_n_142976
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.818 36.317 112.846 36.48 ;
      END
   END FE_OFN13322_n_142976

   PIN FE_OFN13323_n_142975
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.93 36.317 114.958 36.48 ;
      END
   END FE_OFN13323_n_142975

   PIN FE_OFN13325_n_142975
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.018 36.317 108.046 36.48 ;
      END
   END FE_OFN13325_n_142975

   PIN FE_OFN13334_n_142837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.37 36.317 112.398 36.48 ;
      END
   END FE_OFN13334_n_142837

   PIN FE_OFN13341_n_142836
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.506 36.317 123.534 36.48 ;
      END
   END FE_OFN13341_n_142836

   PIN FE_OFN13494_n_111726
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.042 36.317 125.07 36.48 ;
      END
   END FE_OFN13494_n_111726

   PIN FE_OFN13569_n_143090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.714 36.317 113.742 36.48 ;
      END
   END FE_OFN13569_n_143090

   PIN FE_OFN13578_n_143089
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.762 36.317 115.79 36.48 ;
      END
   END FE_OFN13578_n_143089

   PIN FE_OFN13583_n_143088
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.746 36.317 109.774 36.48 ;
      END
   END FE_OFN13583_n_143088

   PIN FE_OFN13590_n_142824
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.57 36.317 115.598 36.48 ;
      END
   END FE_OFN13590_n_142824

   PIN FE_OFN13601_n_142823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.658 36.317 108.686 36.48 ;
      END
   END FE_OFN13601_n_142823

   PIN FE_OFN13734_n_143076
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.922 36.317 103.95 36.48 ;
      END
   END FE_OFN13734_n_143076

   PIN FE_OFN13740_n_143075
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.346 36.317 119.374 36.48 ;
      END
   END FE_OFN13740_n_143075

   PIN FE_OFN13746_n_143074
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.594 36.317 108.622 36.48 ;
      END
   END FE_OFN13746_n_143074

   PIN FE_OFN13753_n_142978
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.642 36.317 110.67 36.48 ;
      END
   END FE_OFN13753_n_142978

   PIN FE_OFN13913_n_111944
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.074 36.317 113.102 36.48 ;
      END
   END FE_OFN13913_n_111944

   PIN FE_OFN14283_n_144177
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.442 36.317 123.47 36.48 ;
      END
   END FE_OFN14283_n_144177

   PIN FE_OFN14445_n_143580
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.53 36.317 100.558 36.48 ;
      END
   END FE_OFN14445_n_143580

   PIN FE_OFN14884_n_590
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 33.522 137.792 33.55 ;
      END
   END FE_OFN14884_n_590

   PIN FE_OFN16411_b_1_4_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.306 36.317 104.334 36.48 ;
      END
   END FE_OFN16411_b_1_4_3

   PIN FE_OFN16414_b_1_4_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.666 36.317 103.694 36.48 ;
      END
   END FE_OFN16414_b_1_4_2

   PIN FE_OFN16657_n_8260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.882 0.163 8.91 ;
      END
   END FE_OFN16657_n_8260

   PIN FE_OFN16659_n_6874
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.378 0.0 19.406 0.163 ;
      END
   END FE_OFN16659_n_6874

   PIN FE_OFN16661_n_8311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.61 0.0 18.638 0.163 ;
      END
   END FE_OFN16661_n_8311

   PIN FE_OFN16665_n_6760
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.586 0.0 17.614 0.163 ;
      END
   END FE_OFN16665_n_6760

   PIN FE_OFN18760_n_142881
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.162 36.317 106.19 36.48 ;
      END
   END FE_OFN18760_n_142881

   PIN FE_OFN18846_n_142838
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.482 36.317 114.51 36.48 ;
      END
   END FE_OFN18846_n_142838

   PIN FE_OFN19317_b_1_0_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.026 36.317 111.054 36.48 ;
      END
   END FE_OFN19317_b_1_0_8

   PIN FE_OFN2291_n_142893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.57 36.317 123.598 36.48 ;
      END
   END FE_OFN2291_n_142893

   PIN FE_OFN2305_n_142891
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.506 36.317 115.534 36.48 ;
      END
   END FE_OFN2305_n_142891

   PIN FE_OFN2501_n_111905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.306 36.317 112.334 36.48 ;
      END
   END FE_OFN2501_n_111905

   PIN FE_OFN2681_n_111726
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.394 36.317 113.422 36.48 ;
      END
   END FE_OFN2681_n_111726

   PIN FE_OFN2697_n_142838
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.874 36.317 109.902 36.48 ;
      END
   END FE_OFN2697_n_142838

   PIN FE_OFN2707_n_142835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.186 36.317 115.214 36.48 ;
      END
   END FE_OFN2707_n_142835

   PIN FE_OFN2766_n_142822
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.538 36.317 111.566 36.48 ;
      END
   END FE_OFN2766_n_142822

   PIN FE_OFN2827_n_142933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.586 36.317 121.614 36.48 ;
      END
   END FE_OFN2827_n_142933

   PIN FE_OFN2887_n_143090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.562 36.317 112.59 36.48 ;
      END
   END FE_OFN2887_n_143090

   PIN FE_OFN3030_n_143115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.906 36.317 97.934 36.48 ;
      END
   END FE_OFN3030_n_143115

   PIN FE_OFN3049_n_143311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.842 36.317 97.87 36.48 ;
      END
   END FE_OFN3049_n_143311

   PIN FE_OFN3057_n_143311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.634 36.317 123.662 36.48 ;
      END
   END FE_OFN3057_n_143311

   PIN FE_OFN558_n_11188
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.106 0.163 5.134 ;
      END
   END FE_OFN558_n_11188

   PIN FE_OFN564_n_8310
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.042 0.163 5.07 ;
      END
   END FE_OFN564_n_8310

   PIN FE_OFN584_n_6873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.338 36.317 12.366 36.48 ;
      END
   END FE_OFN584_n_6873

   PIN FE_OFN934_n_5008
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.722 0.0 12.75 0.163 ;
      END
   END FE_OFN934_n_5008

   PIN b_1_0_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.114 36.317 112.142 36.48 ;
      END
   END b_1_0_0

   PIN b_1_0_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.762 36.317 99.79 36.48 ;
      END
   END b_1_0_1

   PIN b_1_0_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.754 36.317 112.782 36.48 ;
      END
   END b_1_0_10

   PIN b_1_0_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.69 36.317 112.718 36.48 ;
      END
   END b_1_0_4

   PIN b_1_0_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.746 36.317 101.774 36.48 ;
      END
   END b_1_0_6

   PIN b_1_0_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.802 36.317 114.83 36.48 ;
      END
   END b_1_0_9

   PIN b_1_1_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.722 36.317 116.75 36.48 ;
      END
   END b_1_1_10

   PIN b_1_1_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.634 36.317 115.662 36.48 ;
      END
   END b_1_1_11

   PIN b_1_1_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.402 36.317 116.43 36.48 ;
      END
   END b_1_1_12

   PIN b_1_1_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 20.466 137.792 20.494 ;
      END
   END b_1_1_14

   PIN b_1_1_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 112.946 36.317 112.974 36.48 ;
      END
   END b_1_1_2

   PIN b_1_1_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.858 36.317 119.886 36.48 ;
      END
   END b_1_1_3

   PIN b_1_1_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 16.626 137.792 16.654 ;
      END
   END b_1_1_4

   PIN b_1_1_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.378 36.317 123.406 36.48 ;
      END
   END b_1_1_5

   PIN b_1_1_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.786 36.317 124.814 36.48 ;
      END
   END b_1_1_6

   PIN b_1_1_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 131.442 36.317 131.47 36.48 ;
      END
   END b_1_1_7

   PIN b_1_1_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 127.602 36.317 127.63 36.48 ;
      END
   END b_1_1_8

   PIN b_1_1_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.394 36.317 121.422 36.48 ;
      END
   END b_1_1_9

   PIN b_1_3_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 135.282 36.317 135.31 36.48 ;
      END
   END b_1_3_8

   PIN b_1_4_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.378 36.317 115.406 36.48 ;
      END
   END b_1_4_10

   PIN b_1_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.45 36.398 102.478 36.48 ;
      END
   END b_1_4_4

   PIN b_1_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.658 36.317 108.686 36.48 ;
      END
   END b_1_4_5

   PIN b_1_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.73 36.317 103.758 36.48 ;
      END
   END b_1_4_6

   PIN b_1_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.754 36.317 104.782 36.48 ;
      END
   END b_1_4_7

   PIN b_1_4_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.57 36.317 107.598 36.48 ;
      END
   END b_1_4_8

   PIN b_1_4_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.466 36.317 108.494 36.48 ;
      END
   END b_1_4_9

   PIN b_1_9_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.826 36.398 123.854 36.48 ;
      END
   END b_1_9_4

   PIN b_1_9_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 33.586 137.792 33.614 ;
      END
   END b_1_9_6

   PIN b_1_9_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.698 36.317 123.726 36.48 ;
      END
   END b_1_9_9

   PIN delay_add_ln34_unr2_unr9_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.042 0.163 13.07 ;
      END
   END delay_add_ln34_unr2_unr9_stage2_stallmux_z_14_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.314 36.398 3.342 36.48 ;
      END
   END ispd_clk

   PIN mul_4376_72_n_334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.874 36.317 117.902 36.48 ;
      END
   END mul_4376_72_n_334

   PIN mul_4376_72_n_336
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.066 36.317 118.094 36.48 ;
      END
   END mul_4376_72_n_336

   PIN mul_4376_72_n_337
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.682 36.317 117.71 36.48 ;
      END
   END mul_4376_72_n_337

   PIN mul_4376_72_n_766
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.25 36.317 91.278 36.48 ;
      END
   END mul_4376_72_n_766

   PIN mul_4376_72_n_771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.802 36.317 90.83 36.48 ;
      END
   END mul_4376_72_n_771

   PIN mul_4379_72_n_329
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.794 36.317 103.822 36.48 ;
      END
   END mul_4379_72_n_329

   PIN mul_4385_72_n_185
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.282 36.317 103.31 36.48 ;
      END
   END mul_4385_72_n_185

   PIN mul_4385_72_n_218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.266 36.317 97.294 36.48 ;
      END
   END mul_4385_72_n_218

   PIN mul_4385_72_n_288
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.178 36.317 112.206 36.48 ;
      END
   END mul_4385_72_n_288

   PIN mul_4385_72_n_290
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.602 36.317 111.63 36.48 ;
      END
   END mul_4385_72_n_290

   PIN mul_4385_72_n_331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.658 36.317 92.686 36.48 ;
      END
   END mul_4385_72_n_331

   PIN n_10918
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.722 36.317 92.75 36.48 ;
      END
   END n_10918

   PIN n_111893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 28.082 137.792 28.11 ;
      END
   END n_111893

   PIN n_114202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.154 36.317 111.182 36.48 ;
      END
   END n_114202

   PIN n_114322
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.482 36.317 106.51 36.48 ;
      END
   END n_114322

   PIN n_115476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.314 36.317 115.342 36.48 ;
      END
   END n_115476

   PIN n_116062
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.49 36.317 101.518 36.48 ;
      END
   END n_116062

   PIN n_116078
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.554 36.317 109.582 36.48 ;
      END
   END n_116078

   PIN n_116171
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.026 36.317 103.054 36.48 ;
      END
   END n_116171

   PIN n_116178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 119.282 36.317 119.31 36.48 ;
      END
   END n_116178

   PIN n_118837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 109.49 36.317 109.518 36.48 ;
      END
   END n_118837

   PIN n_120395
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.962 36.317 102.99 36.48 ;
      END
   END n_120395

   PIN n_120396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.77 36.317 102.798 36.48 ;
      END
   END n_120396

   PIN n_121024
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.178 36.317 96.206 36.48 ;
      END
   END n_121024

   PIN n_121960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.194 36.317 94.222 36.48 ;
      END
   END n_121960

   PIN n_123542
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.794 36.317 95.822 36.48 ;
      END
   END n_123542

   PIN n_124237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 108.722 36.317 108.75 36.48 ;
      END
   END n_124237

   PIN n_128028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.858 36.317 103.886 36.48 ;
      END
   END n_128028

   PIN n_129300
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.306 36.317 104.334 36.48 ;
      END
   END n_129300

   PIN n_129536
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.05 36.317 104.078 36.48 ;
      END
   END n_129536

   PIN n_140259
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 137.629 33.65 137.792 33.678 ;
      END
   END n_140259

   PIN n_142822
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 116.338 36.317 116.366 36.48 ;
      END
   END n_142822

   PIN n_142894
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.61 36.317 114.638 36.48 ;
      END
   END n_142894

   PIN n_143018
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.194 36.317 118.222 36.48 ;
      END
   END n_143018

   PIN n_143019
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.17 36.317 117.198 36.48 ;
      END
   END n_143019

   PIN n_143638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.322 36.317 118.35 36.48 ;
      END
   END n_143638

   PIN n_14520
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.578 36.317 110.606 36.48 ;
      END
   END n_14520

   PIN n_15473
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.01 36.317 97.038 36.48 ;
      END
   END n_15473

   PIN n_17469
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 121.458 36.317 121.486 36.48 ;
      END
   END n_17469

   PIN n_19194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.09 36.317 71.118 36.48 ;
      END
   END n_19194

   PIN n_276
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.154 36.317 111.182 36.48 ;
      END
   END n_276

   PIN n_31708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.946 36.317 104.974 36.48 ;
      END
   END n_31708

   PIN n_31960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.626 36.317 104.654 36.48 ;
      END
   END n_31960

   PIN n_31969
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.97 36.317 105.998 36.48 ;
      END
   END n_31969

   PIN n_32248
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.21 36.317 108.238 36.48 ;
      END
   END n_32248

   PIN n_32393
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.402 36.317 100.43 36.48 ;
      END
   END n_32393

   PIN n_32609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.786 36.317 116.814 36.48 ;
      END
   END n_32609

   PIN n_33345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.082 36.317 116.11 36.48 ;
      END
   END n_33345

   PIN n_33709
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.226 36.317 106.254 36.48 ;
      END
   END n_33709

   PIN n_35162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.378 36.317 107.406 36.48 ;
      END
   END n_35162

   PIN n_35163
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.314 36.317 107.342 36.48 ;
      END
   END n_35163

   PIN n_36227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.458 36.317 97.486 36.48 ;
      END
   END n_36227

   PIN n_36447
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.586 36.317 97.614 36.48 ;
      END
   END n_36447

   PIN n_36460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.786 36.317 92.814 36.48 ;
      END
   END n_36460

   PIN n_36901
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.57 36.317 123.598 36.48 ;
      END
   END n_36901

   PIN n_37985
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.122 36.317 123.15 36.48 ;
      END
   END n_37985

   PIN n_3815
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.506 36.317 123.534 36.48 ;
      END
   END n_3815

   PIN n_4222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.746 36.317 117.774 36.48 ;
      END
   END n_4222

   PIN n_48966
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.594 36.317 116.622 36.48 ;
      END
   END n_48966

   PIN n_49396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.434 36.317 104.462 36.48 ;
      END
   END n_49396

   PIN n_54005
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.13 36.317 118.158 36.48 ;
      END
   END n_54005

   PIN n_6591
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 127.474 36.317 127.502 36.48 ;
      END
   END n_6591

   PIN n_7713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.698 36.317 115.726 36.48 ;
      END
   END n_7713

   PIN n_7789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.53 36.317 92.558 36.48 ;
      END
   END n_7789

   PIN n_7790
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.386 36.317 110.414 36.48 ;
      END
   END n_7790

   PIN n_8356
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.362 36.317 109.39 36.48 ;
      END
   END n_8356

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 137.792 36.48 ;
      LAYER V1 ;
         RECT 0.0 0.0 137.792 36.48 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 137.792 36.48 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 137.792 36.48 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 137.792 36.48 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 137.792 36.48 ;
      LAYER M1 ;
         RECT 0.0 0.0 137.792 36.48 ;
   END
END h7_mgc_matrix_mult_b

MACRO h6_mgc_matrix_mult_b
   CLASS BLOCK ;
   FOREIGN h6 ;
   ORIGIN 0 0 ;
   SIZE 110.592 BY 116.48 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN15477_n_143101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.266 116.317 105.294 116.48 ;
      END
   END FE_OCPN15477_n_143101

   PIN FE_OCPN15479_n_143101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.706 116.317 102.734 116.48 ;
      END
   END FE_OCPN15479_n_143101

   PIN FE_OFN10194_b_2_8_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.858 116.317 103.886 116.48 ;
      END
   END FE_OFN10194_b_2_8_3

   PIN FE_OFN10197_b_2_8_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.866 116.317 106.894 116.48 ;
      END
   END FE_OFN10197_b_2_8_1

   PIN FE_OFN10200_b_2_8_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.354 116.317 106.382 116.48 ;
      END
   END FE_OFN10200_b_2_8_0

   PIN FE_OFN11317_n_143101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 114.034 110.592 114.062 ;
      END
   END FE_OFN11317_n_143101

   PIN FE_OFN11341_n_142989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.034 116.317 106.062 116.48 ;
      END
   END FE_OFN11341_n_142989

   PIN FE_OFN11351_n_140257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 110.322 110.592 110.35 ;
      END
   END FE_OFN11351_n_140257

   PIN FE_OFN11511_n_143549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 110.258 110.592 110.286 ;
      END
   END FE_OFN11511_n_143549

   PIN FE_OFN11514_n_143549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.458 110.592 113.486 ;
      END
   END FE_OFN11514_n_143549

   PIN FE_OFN11516_n_143549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 107.122 110.592 107.15 ;
      END
   END FE_OFN11516_n_143549

   PIN FE_OFN11593_n_143231
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.394 110.592 113.422 ;
      END
   END FE_OFN11593_n_143231

   PIN FE_OFN11596_n_112428
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 89.458 110.592 89.486 ;
      END
   END FE_OFN11596_n_112428

   PIN FE_OFN11598_n_112428
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 106.482 110.592 106.51 ;
      END
   END FE_OFN11598_n_112428

   PIN FE_OFN11811_n_111876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.162 116.317 106.19 116.48 ;
      END
   END FE_OFN11811_n_111876

   PIN FE_OFN11812_n_111876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.714 110.592 113.742 ;
      END
   END FE_OFN11812_n_111876

   PIN FE_OFN11859_n_143243
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.25 116.317 99.278 116.48 ;
      END
   END FE_OFN11859_n_143243

   PIN FE_OFN11863_n_143230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.386 116.317 102.414 116.48 ;
      END
   END FE_OFN11863_n_143230

   PIN FE_OFN11864_n_143230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.506 116.317 99.534 116.48 ;
      END
   END FE_OFN11864_n_143230

   PIN FE_OFN11886_n_143104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 107.186 110.592 107.214 ;
      END
   END FE_OFN11886_n_143104

   PIN FE_OFN11887_n_143104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.354 116.317 106.382 116.48 ;
      END
   END FE_OFN11887_n_143104

   PIN FE_OFN11888_n_143104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 105.778 110.592 105.806 ;
      END
   END FE_OFN11888_n_143104

   PIN FE_OFN11889_n_143104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 85.618 110.592 85.646 ;
      END
   END FE_OFN11889_n_143104

   PIN FE_OFN11892_n_143103
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.29 116.317 106.318 116.48 ;
      END
   END FE_OFN11892_n_143103

   PIN FE_OFN11893_n_143103
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.33 110.592 113.358 ;
      END
   END FE_OFN11893_n_143103

   PIN FE_OFN11898_n_143062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.986 110.592 112.014 ;
      END
   END FE_OFN11898_n_143062

   PIN FE_OFN11900_n_143062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 115.25 110.592 115.278 ;
      END
   END FE_OFN11900_n_143062

   PIN FE_OFN11901_n_143062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.346 116.317 103.374 116.48 ;
      END
   END FE_OFN11901_n_143062

   PIN FE_OFN11905_n_143061
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 108.722 110.592 108.75 ;
      END
   END FE_OFN11905_n_143061

   PIN FE_OFN11906_n_143061
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 101.234 110.592 101.262 ;
      END
   END FE_OFN11906_n_143061

   PIN FE_OFN11907_n_143060
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 105.202 110.592 105.23 ;
      END
   END FE_OFN11907_n_143060

   PIN FE_OFN11913_n_143060
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.842 116.317 97.87 116.48 ;
      END
   END FE_OFN11913_n_143060

   PIN FE_OFN11920_n_143047
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 85.618 110.592 85.646 ;
      END
   END FE_OFN11920_n_143047

   PIN FE_OFN11921_n_143047
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.29 116.317 106.318 116.48 ;
      END
   END FE_OFN11921_n_143047

   PIN FE_OFN12307_n_111875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 105.906 110.592 105.934 ;
      END
   END FE_OFN12307_n_111875

   PIN FE_OFN12308_n_111875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.354 116.317 98.382 116.48 ;
      END
   END FE_OFN12308_n_111875

   PIN FE_OFN12310_n_111875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.906 116.317 97.934 116.48 ;
      END
   END FE_OFN12310_n_111875

   PIN FE_OFN12312_n_111877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.642 116.317 102.67 116.48 ;
      END
   END FE_OFN12312_n_111877

   PIN FE_OFN12313_n_111877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.13 116.317 102.158 116.48 ;
      END
   END FE_OFN12313_n_111877

   PIN FE_OFN12320_n_112427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.562 110.592 112.59 ;
      END
   END FE_OFN12320_n_112427

   PIN FE_OFN12323_n_112427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.706 116.317 102.734 116.48 ;
      END
   END FE_OFN12323_n_112427

   PIN FE_OFN12325_n_112470
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.818 110.592 112.846 ;
      END
   END FE_OFN12325_n_112470

   PIN FE_OFN12331_n_137473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.97 116.317 105.998 116.48 ;
      END
   END FE_OFN12331_n_137473

   PIN FE_OFN12332_n_137473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.754 110.592 112.782 ;
      END
   END FE_OFN12332_n_137473

   PIN FE_OFN12335_n_137268
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 102.002 110.592 102.03 ;
      END
   END FE_OFN12335_n_137268

   PIN FE_OFN12344_n_142992
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.322 116.317 102.35 116.48 ;
      END
   END FE_OFN12344_n_142992

   PIN FE_OFN12357_n_142922
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 85.554 110.592 85.582 ;
      END
   END FE_OFN12357_n_142922

   PIN FE_OFN12358_n_142922
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 92.594 110.592 92.622 ;
      END
   END FE_OFN12358_n_142922

   PIN FE_OFN12360_n_142922
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 110.386 110.592 110.414 ;
      END
   END FE_OFN12360_n_142922

   PIN FE_OFN12361_n_142922
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.13 116.317 102.158 116.48 ;
      END
   END FE_OFN12361_n_142922

   PIN FE_OFN12365_n_142921
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 101.362 110.592 101.39 ;
      END
   END FE_OFN12365_n_142921

   PIN FE_OFN12366_n_142921
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.51 110.45 110.592 110.478 ;
      END
   END FE_OFN12366_n_142921

   PIN FE_OFN12377_n_142908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.842 116.317 105.87 116.48 ;
      END
   END FE_OFN12377_n_142908

   PIN FE_OFN12378_n_142908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 85.682 110.592 85.71 ;
      END
   END FE_OFN12378_n_142908

   PIN FE_OFN12379_n_142908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.922 110.592 111.95 ;
      END
   END FE_OFN12379_n_142908

   PIN FE_OFN12380_n_142907
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.394 116.317 105.422 116.48 ;
      END
   END FE_OFN12380_n_142907

   PIN FE_OFN12381_n_142907
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 102.066 110.592 102.094 ;
      END
   END FE_OFN12381_n_142907

   PIN FE_OFN12387_n_142906
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.122 110.592 107.15 ;
      END
   END FE_OFN12387_n_142906

   PIN FE_OFN12388_n_142906
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 86.066 110.592 86.094 ;
      END
   END FE_OFN12388_n_142906

   PIN FE_OFN12416_n_143396
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 106.354 110.592 106.382 ;
      END
   END FE_OFN12416_n_143396

   PIN FE_OFN12598_n_111738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 105.97 110.592 105.998 ;
      END
   END FE_OFN12598_n_111738

   PIN FE_OFN12600_n_111738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 109.682 110.592 109.71 ;
      END
   END FE_OFN12600_n_111738

   PIN FE_OFN12601_n_111738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 109.17 110.592 109.198 ;
      END
   END FE_OFN12601_n_111738

   PIN FE_OFN12602_n_111738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.45 116.317 102.478 116.48 ;
      END
   END FE_OFN12602_n_111738

   PIN FE_OFN12607_n_112606
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 110.578 110.592 110.606 ;
      END
   END FE_OFN12607_n_112606

   PIN FE_OFN12608_n_112606
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.066 116.317 102.094 116.48 ;
      END
   END FE_OFN12608_n_112606

   PIN FE_OFN12614_n_112689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.514 116.317 102.542 116.48 ;
      END
   END FE_OFN12614_n_112689

   PIN FE_OFN12615_n_112689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.058 116.317 107.086 116.48 ;
      END
   END FE_OFN12615_n_112689

   PIN FE_OFN12620_n_112690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.794 116.317 103.822 116.48 ;
      END
   END FE_OFN12620_n_112690

   PIN FE_OFN12621_n_112690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.082 110.592 108.11 ;
      END
   END FE_OFN12621_n_112690

   PIN FE_OFN12626_n_143646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.65 116.317 97.678 116.48 ;
      END
   END FE_OFN12626_n_143646

   PIN FE_OFN12653_n_111913
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.842 110.592 113.87 ;
      END
   END FE_OFN12653_n_111913

   PIN FE_OFN12654_n_111913
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.226 116.317 106.254 116.48 ;
      END
   END FE_OFN12654_n_111913

   PIN FE_OFN12655_n_111913
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.69 110.592 112.718 ;
      END
   END FE_OFN12655_n_111913

   PIN FE_OFN13022_n_142949
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 107.442 110.592 107.47 ;
      END
   END FE_OFN13022_n_142949

   PIN FE_OFN13026_n_142948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 99.57 110.592 99.598 ;
      END
   END FE_OFN13026_n_142948

   PIN FE_OFN13027_n_142948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 89.522 110.592 89.55 ;
      END
   END FE_OFN13027_n_142948

   PIN FE_OFN13028_n_142948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.61 116.317 98.638 116.48 ;
      END
   END FE_OFN13028_n_142948

   PIN FE_OFN13554_n_143397
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.626 110.592 104.654 ;
      END
   END FE_OFN13554_n_143397

   PIN FE_OFN13555_n_143397
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 109.106 110.592 109.134 ;
      END
   END FE_OFN13555_n_143397

   PIN FE_OFN13556_n_143397
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 108.53 110.592 108.558 ;
      END
   END FE_OFN13556_n_143397

   PIN FE_OFN15932_n_143241
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.778 116.317 105.806 116.48 ;
      END
   END FE_OFN15932_n_143241

   PIN FE_OFN17143_n_21437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.714 116.317 105.742 116.48 ;
      END
   END FE_OFN17143_n_21437

   PIN FE_OFN17204_n_16278
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.522 116.317 105.55 116.48 ;
      END
   END FE_OFN17204_n_16278

   PIN FE_OFN17229_n_142990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 102.642 110.592 102.67 ;
      END
   END FE_OFN17229_n_142990

   PIN FE_OFN17234_n_142989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 114.866 110.592 114.894 ;
      END
   END FE_OFN17234_n_142989

   PIN FE_OFN18945_n_112470
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.538 110.592 111.566 ;
      END
   END FE_OFN18945_n_112470

   PIN FE_OFN3348_n_14460
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.498 110.592 96.526 ;
      END
   END FE_OFN3348_n_14460

   PIN FE_OFN3417_n_112606
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.338 110.592 108.366 ;
      END
   END FE_OFN3417_n_112606

   PIN FE_OFN3476_n_142921
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.186 116.317 107.214 116.48 ;
      END
   END FE_OFN3476_n_142921

   PIN FE_OFN3535_n_140257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.658 116.317 100.686 116.48 ;
      END
   END FE_OFN3535_n_140257

   PIN FE_OFN3615_n_112427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.802 116.317 106.83 116.48 ;
      END
   END FE_OFN3615_n_112427

   PIN FE_OFN3639_n_143227
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.482 116.317 106.51 116.48 ;
      END
   END FE_OFN3639_n_143227

   PIN FE_OFN3650_n_143231
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.434 110.592 112.462 ;
      END
   END FE_OFN3650_n_143231

   PIN FE_OFN3718_n_143243
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.602 116.317 103.63 116.48 ;
      END
   END FE_OFN3718_n_143243

   PIN FE_OFN3731_n_143397
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 110.962 110.592 110.99 ;
      END
   END FE_OFN3731_n_143397

   PIN FE_OFN3754_n_143549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.57 110.592 107.598 ;
      END
   END FE_OFN3754_n_143549

   PIN FE_OFN3755_n_143549
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.53 110.592 100.558 ;
      END
   END FE_OFN3755_n_143549

   PIN mul_4665_72_n_303
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 93.682 110.592 93.71 ;
      END
   END mul_4665_72_n_303

   PIN mul_4665_72_n_305
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.082 110.592 100.11 ;
      END
   END mul_4665_72_n_305

   PIN mul_4665_72_n_317
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 94.386 110.592 94.414 ;
      END
   END mul_4665_72_n_317

   PIN mul_4665_72_n_318
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 94.45 110.592 94.478 ;
      END
   END mul_4665_72_n_318

   PIN mul_4665_72_n_327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.562 110.592 96.59 ;
      END
   END mul_4665_72_n_327

   PIN mul_4665_72_n_328
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.05 110.592 96.078 ;
      END
   END mul_4665_72_n_328

   PIN mul_4666_72_n_308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 110.962 110.592 110.99 ;
      END
   END mul_4666_72_n_308

   PIN mul_4666_72_n_309
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 108.786 110.592 108.814 ;
      END
   END mul_4666_72_n_309

   PIN mul_4666_72_n_848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.586 116.317 105.614 116.48 ;
      END
   END mul_4666_72_n_848

   PIN mul_4668_72_n_57
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.618 116.317 93.646 116.48 ;
      END
   END mul_4668_72_n_57

   PIN mul_4668_72_n_73
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.554 116.317 93.582 116.48 ;
      END
   END mul_4668_72_n_73

   PIN mul_4668_72_n_767
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.81 116.317 93.838 116.48 ;
      END
   END mul_4668_72_n_767

   PIN mul_4671_72_n_151
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.45 116.317 102.478 116.48 ;
      END
   END mul_4671_72_n_151

   PIN mul_4671_72_n_170
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.194 116.317 102.222 116.48 ;
      END
   END mul_4671_72_n_170

   PIN mul_4671_72_n_225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.186 116.317 91.214 116.48 ;
      END
   END mul_4671_72_n_225

   PIN mul_4671_72_n_251
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.674 116.317 90.702 116.48 ;
      END
   END mul_4671_72_n_251

   PIN mul_4671_72_n_338
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.442 116.317 91.47 116.48 ;
      END
   END mul_4671_72_n_338

   PIN mul_4671_72_n_340
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.57 116.317 91.598 116.48 ;
      END
   END mul_4671_72_n_340

   PIN n_1080
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 91.89 110.592 91.918 ;
      END
   END n_1080

   PIN n_1081
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 91.762 110.592 91.79 ;
      END
   END n_1081

   PIN n_1116
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 91.954 110.592 91.982 ;
      END
   END n_1116

   PIN n_1117
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 92.018 110.592 92.046 ;
      END
   END n_1117

   PIN n_111877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.474 110.592 111.502 ;
      END
   END n_111877

   PIN n_111878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 114.93 110.592 114.958 ;
      END
   END n_111878

   PIN n_11193
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 114.994 110.592 115.022 ;
      END
   END n_11193

   PIN n_112427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.466 110.592 108.494 ;
      END
   END n_112427

   PIN n_112752
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.05 110.592 112.078 ;
      END
   END n_112752

   PIN n_112920
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.442 116.317 107.47 116.48 ;
      END
   END n_112920

   PIN n_113005
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.578 116.317 102.606 116.48 ;
      END
   END n_113005

   PIN n_113236
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.026 116.317 103.054 116.48 ;
      END
   END n_113236

   PIN n_113311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.37 116.317 96.398 116.48 ;
      END
   END n_113311

   PIN n_113414
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.89 116.317 91.918 116.48 ;
      END
   END n_113414

   PIN n_113566
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.994 116.317 99.022 116.48 ;
      END
   END n_113566

   PIN n_113666
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.906 110.592 113.934 ;
      END
   END n_113666

   PIN n_113667
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.162 116.317 106.19 116.48 ;
      END
   END n_113667

   PIN n_113813
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.626 116.317 104.654 116.48 ;
      END
   END n_113813

   PIN n_113885
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.994 116.317 107.022 116.48 ;
      END
   END n_113885

   PIN n_113886
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.178 110.592 112.206 ;
      END
   END n_113886

   PIN n_113889
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.258 116.317 102.286 116.48 ;
      END
   END n_113889

   PIN n_113928
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 103.986 110.592 104.014 ;
      END
   END n_113928

   PIN n_113988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.442 116.317 99.47 116.48 ;
      END
   END n_113988

   PIN n_113989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.458 116.317 105.486 116.48 ;
      END
   END n_113989

   PIN n_114186
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.674 116.317 106.702 116.48 ;
      END
   END n_114186

   PIN n_114247
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.274 110.592 100.302 ;
      END
   END n_114247

   PIN n_114413
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.858 116.317 95.886 116.48 ;
      END
   END n_114413

   PIN n_114864
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 115.058 110.592 115.086 ;
      END
   END n_114864

   PIN n_115329
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.842 116.317 97.87 116.48 ;
      END
   END n_115329

   PIN n_115463
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 105.458 110.592 105.486 ;
      END
   END n_115463

   PIN n_115978
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 94.578 110.592 94.606 ;
      END
   END n_115978

   PIN n_116236
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.034 116.317 106.062 116.48 ;
      END
   END n_116236

   PIN n_118055
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.186 116.317 99.214 116.48 ;
      END
   END n_118055

   PIN n_118083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.61 116.317 106.638 116.48 ;
      END
   END n_118083

   PIN n_118092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.986 116.317 96.014 116.48 ;
      END
   END n_118092

   PIN n_118139
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.05 110.592 104.078 ;
      END
   END n_118139

   PIN n_118170
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.306 116.317 104.334 116.48 ;
      END
   END n_118170

   PIN n_118357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.034 116.317 98.062 116.48 ;
      END
   END n_118357

   PIN n_119785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.138 116.317 105.166 116.48 ;
      END
   END n_119785

   PIN n_119984
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.026 110.592 111.054 ;
      END
   END n_119984

   PIN n_120014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.114 116.317 96.142 116.48 ;
      END
   END n_120014

   PIN n_120034
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.954 116.317 99.982 116.48 ;
      END
   END n_120034

   PIN n_120415
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 102.002 110.592 102.03 ;
      END
   END n_120415

   PIN n_120432
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.794 116.317 95.822 116.48 ;
      END
   END n_120432

   PIN n_120820
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.97 116.317 97.998 116.48 ;
      END
   END n_120820

   PIN n_121838
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.09 110.592 111.118 ;
      END
   END n_121838

   PIN n_121898
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 103.282 110.592 103.31 ;
      END
   END n_121898

   PIN n_122243
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.114 110.592 104.142 ;
      END
   END n_122243

   PIN n_122244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.178 110.592 104.206 ;
      END
   END n_122244

   PIN n_122366
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.674 116.317 98.702 116.48 ;
      END
   END n_122366

   PIN n_122676
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.33 116.317 105.358 116.48 ;
      END
   END n_122676

   PIN n_123562
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.698 116.317 91.726 116.48 ;
      END
   END n_123562

   PIN n_123563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.25 116.317 91.278 116.48 ;
      END
   END n_123563

   PIN n_123583
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.914 110.592 100.942 ;
      END
   END n_123583

   PIN n_123660
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.37 110.592 104.398 ;
      END
   END n_123660

   PIN n_123664
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.434 110.592 104.462 ;
      END
   END n_123664

   PIN n_123911
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.482 116.317 98.51 116.48 ;
      END
   END n_123911

   PIN n_12563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.786 110.592 100.814 ;
      END
   END n_12563

   PIN n_125637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 101.042 110.592 101.07 ;
      END
   END n_125637

   PIN n_126034
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.194 116.317 94.222 116.48 ;
      END
   END n_126034

   PIN n_12651
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 105.586 110.592 105.614 ;
      END
   END n_12651

   PIN n_126615
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.562 110.592 104.59 ;
      END
   END n_126615

   PIN n_126616
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 105.266 110.592 105.294 ;
      END
   END n_126616

   PIN n_126766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.738 116.317 90.766 116.48 ;
      END
   END n_126766

   PIN n_127005
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.234 116.317 93.262 116.48 ;
      END
   END n_127005

   PIN n_128115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.778 116.317 97.806 116.48 ;
      END
   END n_128115

   PIN n_129077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.29 116.317 90.318 116.48 ;
      END
   END n_129077

   PIN n_129225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.914 116.317 92.942 116.48 ;
      END
   END n_129225

   PIN n_129226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.042 116.317 93.07 116.48 ;
      END
   END n_129226

   PIN n_129237
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 115.122 110.592 115.15 ;
      END
   END n_129237

   PIN n_130207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 97.65 110.592 97.678 ;
      END
   END n_130207

   PIN n_130208
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 97.714 110.592 97.742 ;
      END
   END n_130208

   PIN n_131285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 93.81 110.592 93.838 ;
      END
   END n_131285

   PIN n_131287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.658 110.592 100.686 ;
      END
   END n_131287

   PIN n_131292
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.954 116.317 91.982 116.48 ;
      END
   END n_131292

   PIN n_131450
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.394 116.317 89.422 116.48 ;
      END
   END n_131450

   PIN n_133179
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 97.074 110.592 97.102 ;
      END
   END n_133179

   PIN n_133200
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 102.066 110.592 102.094 ;
      END
   END n_133200

   PIN n_133250
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.226 116.317 90.254 116.48 ;
      END
   END n_133250

   PIN n_133423
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.73 116.317 95.758 116.48 ;
      END
   END n_133423

   PIN n_133476
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.338 110.592 100.366 ;
      END
   END n_133476

   PIN n_134206
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.434 110.592 96.462 ;
      END
   END n_134206

   PIN n_134263
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.242 116.317 88.27 116.48 ;
      END
   END n_134263

   PIN n_135022
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.306 116.317 88.334 116.48 ;
      END
   END n_135022

   PIN n_13640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 78.066 110.592 78.094 ;
      END
   END n_13640

   PIN n_142908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.906 116.317 105.934 116.48 ;
      END
   END n_142908

   PIN n_142909
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.138 110.592 113.166 ;
      END
   END n_142909

   PIN n_142949
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.274 110.592 108.302 ;
      END
   END n_142949

   PIN n_142990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 105.842 110.592 105.87 ;
      END
   END n_142990

   PIN n_143047
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 106.482 110.592 106.51 ;
      END
   END n_143047

   PIN n_143103
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 101.426 110.592 101.454 ;
      END
   END n_143103

   PIN n_143105
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.122 116.317 107.15 116.48 ;
      END
   END n_143105

   PIN n_143227
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.51 111.346 110.592 111.374 ;
      END
   END n_143227

   PIN n_143230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 97.074 110.592 97.102 ;
      END
   END n_143230

   PIN n_143399
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 109.81 110.592 109.838 ;
      END
   END n_143399

   PIN n_144318
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 62.642 110.592 62.67 ;
      END
   END n_144318

   PIN n_144319
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.986 116.317 104.014 116.48 ;
      END
   END n_144319

   PIN n_14458
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 98.802 110.592 98.83 ;
      END
   END n_14458

   PIN n_14498
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.626 110.592 96.654 ;
      END
   END n_14498

   PIN n_14596
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 99.442 110.592 99.47 ;
      END
   END n_14596

   PIN n_14610
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 89.33 110.592 89.358 ;
      END
   END n_14610

   PIN n_15054
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 81.778 110.592 81.806 ;
      END
   END n_15054

   PIN n_16295
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 101.49 110.592 101.518 ;
      END
   END n_16295

   PIN n_16449
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 93.746 110.592 93.774 ;
      END
   END n_16449

   PIN n_16450
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 94.642 110.592 94.67 ;
      END
   END n_16450

   PIN n_16451
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 94.514 110.592 94.542 ;
      END
   END n_16451

   PIN n_17519
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 89.202 110.592 89.23 ;
      END
   END n_17519

   PIN n_17521
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 89.842 110.592 89.87 ;
      END
   END n_17521

   PIN n_18074
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 86.002 110.592 86.03 ;
      END
   END n_18074

   PIN n_18268
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 93.042 110.592 93.07 ;
      END
   END n_18268

   PIN n_18269
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 93.234 110.592 93.262 ;
      END
   END n_18269

   PIN n_18270
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 93.298 110.592 93.326 ;
      END
   END n_18270

   PIN n_18271
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 89.906 110.592 89.934 ;
      END
   END n_18271

   PIN n_20858
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.482 116.317 106.51 116.48 ;
      END
   END n_20858

   PIN n_20869
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.738 116.317 106.766 116.48 ;
      END
   END n_20869

   PIN n_2993
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.498 110.592 104.526 ;
      END
   END n_2993

   PIN n_3080
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.074 110.592 113.102 ;
      END
   END n_3080

   PIN n_3081
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.946 110.592 112.974 ;
      END
   END n_3081

   PIN n_32762
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.194 116.317 102.222 116.48 ;
      END
   END n_32762

   PIN n_33403
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.01 110.592 113.038 ;
      END
   END n_33403

   PIN n_33960
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.85 116.317 100.878 116.48 ;
      END
   END n_33960

   PIN n_34015
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.106 116.317 101.134 116.48 ;
      END
   END n_34015

   PIN n_34242
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.682 116.317 101.71 116.48 ;
      END
   END n_34242

   PIN n_3519
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 108.018 110.592 108.046 ;
      END
   END n_3519

   PIN n_3543
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.154 110.592 111.182 ;
      END
   END n_3543

   PIN n_3620
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.73 110.592 111.758 ;
      END
   END n_3620

   PIN n_372
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 97.138 110.592 97.166 ;
      END
   END n_372

   PIN n_3728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.57 116.317 107.598 116.48 ;
      END
   END n_3728

   PIN n_3823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.778 110.592 113.806 ;
      END
   END n_3823

   PIN n_3824
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.65 110.592 113.678 ;
      END
   END n_3824

   PIN n_3915
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.242 110.592 96.27 ;
      END
   END n_3915

   PIN n_39274
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.634 110.592 107.662 ;
      END
   END n_39274

   PIN n_5066
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.21 110.592 108.238 ;
      END
   END n_5066

   PIN n_5085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.866 116.317 106.894 116.48 ;
      END
   END n_5085

   PIN n_5164
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 110.45 110.592 110.478 ;
      END
   END n_5164

   PIN n_5958
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 81.97 110.592 81.998 ;
      END
   END n_5958

   PIN n_6550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 108.082 110.592 108.11 ;
      END
   END n_6550

   PIN n_6837
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.954 116.317 99.982 116.48 ;
      END
   END n_6837

   PIN n_6937
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 58.802 110.592 58.83 ;
      END
   END n_6937

   PIN n_8246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.794 110.592 111.822 ;
      END
   END n_8246

   PIN n_8247
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 58.866 110.592 58.894 ;
      END
   END n_8247

   PIN n_8251
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 106.226 110.592 106.254 ;
      END
   END n_8251

   PIN n_8256
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.402 110.592 108.43 ;
      END
   END n_8256

   PIN n_8312
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.146 110.592 108.174 ;
      END
   END n_8312

   PIN n_8343
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 62.706 110.592 62.734 ;
      END
   END n_8343

   PIN n_8481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 84.722 110.592 84.75 ;
      END
   END n_8481

   PIN n_8788
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.658 110.592 108.686 ;
      END
   END n_8788

   PIN n_8789
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 109.746 110.592 109.774 ;
      END
   END n_8789

   PIN n_976
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 93.106 110.592 93.134 ;
      END
   END n_976

   PIN FE_OFN10190_b_2_9_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.226 116.317 106.254 116.48 ;
      END
   END FE_OFN10190_b_2_9_2

   PIN FE_OFN10235_b_2_5_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.322 116.317 102.35 116.48 ;
      END
   END FE_OFN10235_b_2_5_6

   PIN FE_OFN10237_b_2_5_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.978 116.317 101.006 116.48 ;
      END
   END FE_OFN10237_b_2_5_5

   PIN FE_OFN10240_b_2_5_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.722 116.317 100.75 116.48 ;
      END
   END FE_OFN10240_b_2_5_4

   PIN FE_OFN10242_b_2_5_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.786 116.317 100.814 116.48 ;
      END
   END FE_OFN10242_b_2_5_3

   PIN FE_OFN10244_b_2_5_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.938 116.317 101.966 116.48 ;
      END
   END FE_OFN10244_b_2_5_2

   PIN FE_OFN10247_b_2_5_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.674 116.317 106.702 116.48 ;
      END
   END FE_OFN10247_b_2_5_1

   PIN FE_OFN10252_b_2_5_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.498 110.592 112.526 ;
      END
   END FE_OFN10252_b_2_5_0

   PIN FE_OFN10253_b_2_5_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.57 116.317 99.598 116.48 ;
      END
   END FE_OFN10253_b_2_5_0

   PIN FE_OFN10286_b_2_3_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.602 110.592 111.63 ;
      END
   END FE_OFN10286_b_2_3_1

   PIN FE_OFN10288_b_2_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 108.402 110.592 108.43 ;
      END
   END FE_OFN10288_b_2_3_0

   PIN FE_OFN10295_b_2_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 97.01 110.592 97.038 ;
      END
   END FE_OFN10295_b_2_2_2

   PIN FE_OFN10302_b_2_1_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 81.906 110.592 81.934 ;
      END
   END FE_OFN10302_b_2_1_6

   PIN FE_OFN10304_b_2_1_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 82.034 110.592 82.062 ;
      END
   END FE_OFN10304_b_2_1_5

   PIN FE_OFN10306_b_2_1_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 86.13 110.592 86.158 ;
      END
   END FE_OFN10306_b_2_1_4

   PIN FE_OFN10308_b_2_1_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 90.162 110.592 90.19 ;
      END
   END FE_OFN10308_b_2_1_3

   PIN FE_OFN10312_b_2_1_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 91.826 110.592 91.854 ;
      END
   END FE_OFN10312_b_2_1_1

   PIN FE_OFN10314_b_2_1_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 92.402 110.592 92.43 ;
      END
   END FE_OFN10314_b_2_1_0

   PIN FE_OFN11316_n_143101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 114.802 110.592 114.83 ;
      END
   END FE_OFN11316_n_143101

   PIN FE_OFN11338_n_143645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 101.106 110.592 101.134 ;
      END
   END FE_OFN11338_n_143645

   PIN FE_OFN11339_n_142989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.33 116.317 105.358 116.48 ;
      END
   END FE_OFN11339_n_142989

   PIN FE_OFN11365_n_112550
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.378 116.317 107.406 116.48 ;
      END
   END FE_OFN11365_n_112550

   PIN FE_OFN11397_n_140245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.954 110.592 107.982 ;
      END
   END FE_OFN11397_n_140245

   PIN FE_OFN11428_n_142905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.586 116.317 105.614 116.48 ;
      END
   END FE_OFN11428_n_142905

   PIN FE_OFN11429_n_142905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 112.242 110.592 112.27 ;
      END
   END FE_OFN11429_n_142905

   PIN FE_OFN11435_n_142919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 113.138 110.592 113.166 ;
      END
   END FE_OFN11435_n_142919

   PIN FE_OFN11706_n_142947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.394 116.317 97.422 116.48 ;
      END
   END FE_OFN11706_n_142947

   PIN FE_OFN11857_n_143243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.21 110.592 100.238 ;
      END
   END FE_OFN11857_n_143243

   PIN FE_OFN11871_n_143229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 115.378 110.592 115.406 ;
      END
   END FE_OFN11871_n_143229

   PIN FE_OFN11875_n_143227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 97.01 110.592 97.038 ;
      END
   END FE_OFN11875_n_143227

   PIN FE_OFN11876_n_143227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.51 92.21 110.592 92.238 ;
      END
   END FE_OFN11876_n_143227

   PIN FE_OFN11896_n_143102
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 113.074 110.592 113.102 ;
      END
   END FE_OFN11896_n_143102

   PIN FE_OFN11903_n_143061
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.202 110.592 113.23 ;
      END
   END FE_OFN11903_n_143061

   PIN FE_OFN11917_n_143048
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 86.002 110.592 86.03 ;
      END
   END FE_OFN11917_n_143048

   PIN FE_OFN11923_n_143047
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.898 116.317 102.926 116.48 ;
      END
   END FE_OFN11923_n_143047

   PIN FE_OFN12333_n_137473
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 111.602 110.592 111.63 ;
      END
   END FE_OFN12333_n_137473

   PIN FE_OFN12336_n_137268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.51 90.802 110.592 90.83 ;
      END
   END FE_OFN12336_n_137268

   PIN FE_OFN12343_n_142992
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 114.738 110.592 114.766 ;
      END
   END FE_OFN12343_n_142992

   PIN FE_OFN12348_n_142991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 113.01 110.592 113.038 ;
      END
   END FE_OFN12348_n_142991

   PIN FE_OFN12349_n_142991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 110.13 110.592 110.158 ;
      END
   END FE_OFN12349_n_142991

   PIN FE_OFN12350_n_142991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 91.122 110.592 91.15 ;
      END
   END FE_OFN12350_n_142991

   PIN FE_OFN12369_n_142920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 115.314 110.592 115.342 ;
      END
   END FE_OFN12369_n_142920

   PIN FE_OFN12371_n_142920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 90.098 110.592 90.126 ;
      END
   END FE_OFN12371_n_142920

   PIN FE_OFN12374_n_142920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 110.066 110.592 110.094 ;
      END
   END FE_OFN12374_n_142920

   PIN FE_OFN12384_n_142907
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 85.362 110.592 85.39 ;
      END
   END FE_OFN12384_n_142907

   PIN FE_OFN12385_n_142906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 106.29 110.592 106.318 ;
      END
   END FE_OFN12385_n_142906

   PIN FE_OFN12399_n_620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 95.666 110.592 95.694 ;
      END
   END FE_OFN12399_n_620

   PIN FE_OFN12401_n_694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.51 112.882 110.592 112.91 ;
      END
   END FE_OFN12401_n_694

   PIN FE_OFN12595_n_111737
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 108.594 110.592 108.622 ;
      END
   END FE_OFN12595_n_111737

   PIN FE_OFN12612_n_112608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.51 99.442 110.592 99.47 ;
      END
   END FE_OFN12612_n_112608

   PIN FE_OFN12625_n_143646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 89.266 110.592 89.294 ;
      END
   END FE_OFN12625_n_143646

   PIN FE_OFN13015_n_142950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 96.69 110.592 96.718 ;
      END
   END FE_OFN13015_n_142950

   PIN FE_OFN13019_n_142949
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 101.298 110.592 101.326 ;
      END
   END FE_OFN13019_n_142949

   PIN FE_OFN13021_n_142949
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 93.17 110.592 93.198 ;
      END
   END FE_OFN13021_n_142949

   PIN FE_OFN14267_n_140244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 93.234 110.592 93.262 ;
      END
   END FE_OFN14267_n_140244

   PIN FE_OFN14364_n_372
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 89.202 110.592 89.23 ;
      END
   END FE_OFN14364_n_372

   PIN FE_OFN14471_n_143059
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.674 116.317 98.702 116.48 ;
      END
   END FE_OFN14471_n_143059

   PIN FE_OFN14925_n_142989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 90.482 110.592 90.51 ;
      END
   END FE_OFN14925_n_142989

   PIN FE_OFN14959_n_142989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.53 116.317 100.558 116.48 ;
      END
   END FE_OFN14959_n_142989

   PIN FE_OFN15931_n_143241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 114.674 110.592 114.702 ;
      END
   END FE_OFN15931_n_143241

   PIN FE_OFN17142_n_21437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 114.61 110.592 114.638 ;
      END
   END FE_OFN17142_n_21437

   PIN FE_OFN17225_n_140257
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.994 116.317 107.022 116.48 ;
      END
   END FE_OFN17225_n_140257

   PIN FE_OFN17260_n_140245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 105.714 110.592 105.742 ;
      END
   END FE_OFN17260_n_140245

   PIN FE_OFN17262_n_140245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.57 116.317 99.598 116.48 ;
      END
   END FE_OFN17262_n_140245

   PIN FE_OFN18609_b_2_2_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 95.858 110.592 95.886 ;
      END
   END FE_OFN18609_b_2_2_0

   PIN FE_OFN18613_b_2_1_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 92.402 110.592 92.43 ;
      END
   END FE_OFN18613_b_2_1_2

   PIN FE_OFN19151_n_140244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 103.922 110.592 103.95 ;
      END
   END FE_OFN19151_n_140244

   PIN FE_OFN19152_n_890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.242 110.592 112.27 ;
      END
   END FE_OFN19152_n_890

   PIN FE_OFN2212_n_19616
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.458 116.317 105.486 116.48 ;
      END
   END FE_OFN2212_n_19616

   PIN FE_OFN2267_n_19602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.61 116.317 106.638 116.48 ;
      END
   END FE_OFN2267_n_19602

   PIN FE_OFN3491_n_142919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.914 116.317 100.942 116.48 ;
      END
   END FE_OFN3491_n_142919

   PIN FE_OFN3531_n_372
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 96.626 110.592 96.654 ;
      END
   END FE_OFN3531_n_372

   PIN FE_OFN3632_n_143045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.466 110.592 100.494 ;
      END
   END FE_OFN3632_n_143045

   PIN FE_OFN3654_n_112550
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.074 116.317 97.102 116.48 ;
      END
   END FE_OFN3654_n_112550

   PIN FE_OFN3723_n_143241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 110.578 110.592 110.606 ;
      END
   END FE_OFN3723_n_143241

   PIN FE_OFN3746_n_143551
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.018 116.317 100.046 116.48 ;
      END
   END FE_OFN3746_n_143551

   PIN FE_OFN3767_n_143645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 98.162 110.592 98.19 ;
      END
   END FE_OFN3767_n_143645

   PIN b_2_2_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.506 110.592 107.534 ;
      END
   END b_2_2_10

   PIN b_2_2_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.058 0.0 107.086 0.163 ;
      END
   END b_2_2_11

   PIN b_2_2_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.85 110.592 100.878 ;
      END
   END b_2_2_12

   PIN b_2_2_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.906 0.0 105.934 0.163 ;
      END
   END b_2_2_13

   PIN b_2_2_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.906 0.0 105.934 0.163 ;
      END
   END b_2_2_14

   PIN b_2_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 98.29 110.592 98.318 ;
      END
   END b_2_2_3

   PIN b_2_2_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 66.546 110.592 66.574 ;
      END
   END b_2_2_5

   PIN b_2_2_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.978 110.592 101.006 ;
      END
   END b_2_2_6

   PIN b_2_2_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 97.586 110.592 97.614 ;
      END
   END b_2_2_7

   PIN b_2_2_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 98.802 110.592 98.83 ;
      END
   END b_2_2_8

   PIN b_2_2_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 95.09 110.592 95.118 ;
      END
   END b_2_2_9

   PIN b_2_3_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 108.466 110.592 108.494 ;
      END
   END b_2_3_2

   PIN b_2_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 105.842 110.592 105.87 ;
      END
   END b_2_3_3

   PIN b_2_3_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.306 110.592 112.334 ;
      END
   END b_2_3_4

   PIN b_2_3_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.762 110.592 107.79 ;
      END
   END b_2_3_5

   PIN b_2_3_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.098 116.317 106.126 116.48 ;
      END
   END b_2_3_9

   PIN b_2_5_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 114.098 110.592 114.126 ;
      END
   END b_2_5_12

   PIN b_2_5_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 95.794 110.592 95.822 ;
      END
   END b_2_5_8

   PIN b_2_8_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.354 116.317 98.382 116.48 ;
      END
   END b_2_8_0

   PIN b_2_8_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.61 116.317 98.638 116.48 ;
      END
   END b_2_8_1

   PIN b_2_8_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 97.202 110.592 97.23 ;
      END
   END b_2_8_10

   PIN b_2_8_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 96.05 116.317 96.078 116.48 ;
      END
   END b_2_8_11

   PIN b_2_8_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.13 0.0 102.158 0.163 ;
      END
   END b_2_8_12

   PIN b_2_8_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.13 0.0 102.158 0.163 ;
      END
   END b_2_8_13

   PIN b_2_8_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.066 0.0 102.094 0.163 ;
      END
   END b_2_8_14

   PIN b_2_8_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.834 116.317 102.862 116.48 ;
      END
   END b_2_8_2

   PIN b_2_8_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.922 116.317 95.95 116.48 ;
      END
   END b_2_8_3

   PIN b_2_8_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.402 110.592 100.43 ;
      END
   END b_2_8_4

   PIN b_2_8_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.474 116.398 103.502 116.48 ;
      END
   END b_2_8_5

   PIN b_2_8_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.098 116.317 98.126 116.48 ;
      END
   END b_2_8_6

   PIN b_2_8_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.77 116.317 102.798 116.48 ;
      END
   END b_2_8_7

   PIN b_2_8_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.586 116.317 97.614 116.48 ;
      END
   END b_2_8_8

   PIN b_2_8_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.002 0.0 102.03 0.163 ;
      END
   END b_2_8_9

   PIN b_2_9_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.418 116.317 106.446 116.48 ;
      END
   END b_2_9_10

   PIN b_2_9_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.51 96.882 110.592 96.91 ;
      END
   END b_2_9_3

   PIN b_2_9_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.51 114.418 110.592 114.446 ;
      END
   END b_2_9_4

   PIN b_2_9_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 114.29 110.592 114.318 ;
      END
   END b_2_9_6

   PIN b_2_9_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 97.522 110.592 97.55 ;
      END
   END b_2_9_7

   PIN b_2_9_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 111.666 110.592 111.694 ;
      END
   END b_2_9_9

   PIN mul_4665_72_n_306
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.146 110.592 100.174 ;
      END
   END mul_4665_72_n_306

   PIN mul_4665_72_n_326
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.37 110.592 96.398 ;
      END
   END mul_4665_72_n_326

   PIN mul_4665_72_n_332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 101.17 110.592 101.198 ;
      END
   END mul_4665_72_n_332

   PIN mul_4665_72_n_334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.946 110.592 96.974 ;
      END
   END mul_4665_72_n_334

   PIN mul_4666_72_n_73
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.906 116.317 105.934 116.48 ;
      END
   END mul_4666_72_n_73

   PIN mul_4671_72_n_319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.546 116.317 98.574 116.48 ;
      END
   END mul_4671_72_n_319

   PIN n_1001
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 93.17 110.592 93.198 ;
      END
   END n_1001

   PIN n_10204
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 81.842 110.592 81.87 ;
      END
   END n_10204

   PIN n_10206
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 85.49 110.592 85.518 ;
      END
   END n_10206

   PIN n_1038
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 92.082 110.592 92.11 ;
      END
   END n_1038

   PIN n_10399
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 94.962 110.592 94.99 ;
      END
   END n_10399

   PIN n_10464
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 95.602 110.592 95.63 ;
      END
   END n_10464

   PIN n_1075
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 88.37 110.592 88.398 ;
      END
   END n_1075

   PIN n_1099
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 88.178 110.592 88.206 ;
      END
   END n_1099

   PIN n_111913
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 110.514 110.592 110.542 ;
      END
   END n_111913

   PIN n_112428
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 98.226 110.592 98.254 ;
      END
   END n_112428

   PIN n_112607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.51 106.098 110.592 106.126 ;
      END
   END n_112607

   PIN n_112689
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 108.85 110.592 108.878 ;
      END
   END n_112689

   PIN n_113107
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.714 116.317 97.742 116.48 ;
      END
   END n_113107

   PIN n_113124
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.69 116.317 104.718 116.48 ;
      END
   END n_113124

   PIN n_113125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.37 116.317 104.398 116.48 ;
      END
   END n_113125

   PIN n_113149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 109.49 110.592 109.518 ;
      END
   END n_113149

   PIN n_113413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.594 110.592 100.622 ;
      END
   END n_113413

   PIN n_113987
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.506 116.317 99.534 116.48 ;
      END
   END n_113987

   PIN n_114013
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.258 116.317 102.286 116.48 ;
      END
   END n_114013

   PIN n_114266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 106.29 110.592 106.318 ;
      END
   END n_114266

   PIN n_115328
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.906 116.317 97.934 116.48 ;
      END
   END n_115328

   PIN n_115332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.586 116.317 97.614 116.48 ;
      END
   END n_115332

   PIN n_116920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 105.65 110.592 105.678 ;
      END
   END n_116920

   PIN n_118138
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.034 116.317 90.062 116.48 ;
      END
   END n_118138

   PIN n_118140
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 103.602 110.592 103.63 ;
      END
   END n_118140

   PIN n_119676
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 100.722 110.592 100.75 ;
      END
   END n_119676

   PIN n_119760
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 105.33 110.592 105.358 ;
      END
   END n_119760

   PIN n_119922
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.498 116.317 96.526 116.48 ;
      END
   END n_119922

   PIN n_119923
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.714 116.317 97.742 116.48 ;
      END
   END n_119923

   PIN n_121953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.322 116.317 94.35 116.48 ;
      END
   END n_121953

   PIN n_122725
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.666 116.317 95.694 116.48 ;
      END
   END n_122725

   PIN n_12357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 115.186 110.592 115.214 ;
      END
   END n_12357

   PIN n_123790
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.802 116.317 106.83 116.48 ;
      END
   END n_123790

   PIN n_123797
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 104.306 110.592 104.334 ;
      END
   END n_123797

   PIN n_123901
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.93 116.317 90.958 116.48 ;
      END
   END n_123901

   PIN n_124234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.258 116.317 94.286 116.48 ;
      END
   END n_124234

   PIN n_124239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.154 116.317 95.182 116.48 ;
      END
   END n_124239

   PIN n_124242
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.282 116.317 95.31 116.48 ;
      END
   END n_124242

   PIN n_124243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.77 116.317 94.798 116.48 ;
      END
   END n_124243

   PIN n_124266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.586 110.592 113.614 ;
      END
   END n_124266

   PIN n_124799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.842 116.317 89.87 116.48 ;
      END
   END n_124799

   PIN n_125460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 113.522 110.592 113.55 ;
      END
   END n_125460

   PIN n_126110
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.13 116.317 94.158 116.48 ;
      END
   END n_126110

   PIN n_127002
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.106 116.317 93.134 116.48 ;
      END
   END n_127002

   PIN n_127003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.298 116.317 93.326 116.48 ;
      END
   END n_127003

   PIN n_127585
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 112.882 110.592 112.91 ;
      END
   END n_127585

   PIN n_129236
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 114.546 110.592 114.574 ;
      END
   END n_129236

   PIN n_131286
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 101.362 110.592 101.39 ;
      END
   END n_131286

   PIN n_132107
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 94.322 110.592 94.35 ;
      END
   END n_132107

   PIN n_133429
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.826 116.317 91.854 116.48 ;
      END
   END n_133429

   PIN n_134203
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 95.73 110.592 95.758 ;
      END
   END n_134203

   PIN n_134205
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.306 110.592 96.334 ;
      END
   END n_134205

   PIN n_134261
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.586 116.317 89.614 116.48 ;
      END
   END n_134261

   PIN n_134791
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.37 116.317 88.398 116.48 ;
      END
   END n_134791

   PIN n_142907
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 114.226 110.592 114.254 ;
      END
   END n_142907

   PIN n_142993
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 104.946 116.317 104.974 116.48 ;
      END
   END n_142993

   PIN n_143060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 109.042 110.592 109.07 ;
      END
   END n_143060

   PIN n_143063
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.842 116.317 105.87 116.48 ;
      END
   END n_143063

   PIN n_143101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.97 116.317 105.998 116.48 ;
      END
   END n_143101

   PIN n_143231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 106.418 116.317 106.446 116.48 ;
      END
   END n_143231

   PIN n_143396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.442 110.592 107.47 ;
      END
   END n_143396

   PIN n_143549
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.266 116.317 105.294 116.48 ;
      END
   END n_143549

   PIN n_143646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 96.882 110.592 96.91 ;
      END
   END n_143646

   PIN n_14374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.314 116.317 107.342 116.48 ;
      END
   END n_14374

   PIN n_16043
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.546 116.317 106.574 116.48 ;
      END
   END n_16043

   PIN n_1610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 86.194 110.592 86.222 ;
      END
   END n_1610

   PIN n_16278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 114.162 110.592 114.19 ;
      END
   END n_16278

   PIN n_16346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 110.194 110.592 110.222 ;
      END
   END n_16346

   PIN n_3153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 74.226 110.592 74.254 ;
      END
   END n_3153

   PIN n_3207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.89 110.592 107.918 ;
      END
   END n_3207

   PIN n_3208
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.826 110.592 107.854 ;
      END
   END n_3208

   PIN n_32761
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.554 116.317 101.582 116.48 ;
      END
   END n_32761

   PIN n_3404
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 110.429 94.642 110.592 94.67 ;
      END
   END n_3404

   PIN n_3447
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 74.162 110.592 74.19 ;
      END
   END n_3447

   PIN n_3489
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.378 110.592 107.406 ;
      END
   END n_3489

   PIN n_3490
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.314 110.592 107.342 ;
      END
   END n_3490

   PIN n_3813
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.25 110.592 107.278 ;
      END
   END n_3813

   PIN n_3814
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 107.186 110.592 107.214 ;
      END
   END n_3814

   PIN n_3916
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 94.962 110.592 94.99 ;
      END
   END n_3916

   PIN n_3946
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 95.026 110.592 95.054 ;
      END
   END n_3946

   PIN n_5163
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 110.429 110.322 110.592 110.35 ;
      END
   END n_5163

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 110.592 116.48 ;
      LAYER V1 ;
         RECT 0.0 0.0 110.592 116.48 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 110.592 116.48 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 110.592 116.48 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 110.592 116.48 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 110.592 116.48 ;
      LAYER M1 ;
         RECT 0.0 0.0 110.592 116.48 ;
   END
END h6_mgc_matrix_mult_b

MACRO h2_mgc_matrix_mult_b
   CLASS BLOCK ;
   FOREIGN h2 ;
   ORIGIN 0 0 ;
   SIZE 249.792 BY 117.76 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN10016_b_4_4_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.314 0.0 51.342 0.163 ;
      END
   END FE_OFN10016_b_4_4_7

   PIN FE_OFN10107_b_4_2_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.402 0.0 60.43 0.163 ;
      END
   END FE_OFN10107_b_4_2_1

   PIN FE_OFN11689_n_140213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 15.474 249.792 15.502 ;
      END
   END FE_OFN11689_n_140213

   PIN FE_OFN11938_n_142850
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.05 0.0 96.078 0.163 ;
      END
   END FE_OFN11938_n_142850

   PIN FE_OFN12338_n_41013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.626 249.792 48.654 ;
      END
   END FE_OFN12338_n_41013

   PIN FE_OFN12341_n_41013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.898 249.792 30.926 ;
      END
   END FE_OFN12341_n_41013

   PIN FE_OFN12622_n_143670
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.074 249.792 41.102 ;
      END
   END FE_OFN12622_n_143670

   PIN FE_OFN12767_n_41734
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 53.362 249.792 53.39 ;
      END
   END FE_OFN12767_n_41734

   PIN FE_OFN12972_n_41962
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 38.258 249.792 38.286 ;
      END
   END FE_OFN12972_n_41962

   PIN FE_OFN13039_n_40828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.77 249.792 22.798 ;
      END
   END FE_OFN13039_n_40828

   PIN FE_OFN13195_n_137475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 18.482 249.792 18.51 ;
      END
   END FE_OFN13195_n_137475

   PIN FE_OFN13196_n_137475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 64.946 249.792 64.974 ;
      END
   END FE_OFN13196_n_137475

   PIN FE_OFN13200_n_137235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 8.178 249.792 8.206 ;
      END
   END FE_OFN13200_n_137235

   PIN FE_OFN13211_n_143630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 8.242 249.792 8.27 ;
      END
   END FE_OFN13211_n_143630

   PIN FE_OFN13228_n_143481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.65 249.792 57.678 ;
      END
   END FE_OFN13228_n_143481

   PIN FE_OFN13229_n_143481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 69.042 249.792 69.07 ;
      END
   END FE_OFN13229_n_143481

   PIN FE_OFN13244_n_41374
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 53.81 249.792 53.838 ;
      END
   END FE_OFN13244_n_41374

   PIN FE_OFN13247_n_143370
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.93 249.792 26.958 ;
      END
   END FE_OFN13247_n_143370

   PIN FE_OFN13354_n_41014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.09 249.792 55.118 ;
      END
   END FE_OFN13354_n_41014

   PIN FE_OFN13387_n_41612
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 45.938 249.792 45.966 ;
      END
   END FE_OFN13387_n_41612

   PIN FE_OFN13390_n_41612
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.258 249.792 30.286 ;
      END
   END FE_OFN13390_n_41612

   PIN FE_OFN13420_n_41709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 61.106 249.792 61.134 ;
      END
   END FE_OFN13420_n_41709

   PIN FE_OFN13421_n_41709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.834 249.792 22.862 ;
      END
   END FE_OFN13421_n_41709

   PIN FE_OFN13527_n_137233
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.026 249.792 15.054 ;
      END
   END FE_OFN13527_n_137233

   PIN FE_OFN13530_n_137233
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.674 249.792 26.702 ;
      END
   END FE_OFN13530_n_137233

   PIN FE_OFN13619_n_41963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.898 249.792 22.926 ;
      END
   END FE_OFN13619_n_41963

   PIN FE_OFN13620_n_41963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.946 249.792 80.974 ;
      END
   END FE_OFN13620_n_41963

   PIN FE_OFN13621_n_41963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 4.082 249.792 4.11 ;
      END
   END FE_OFN13621_n_41963

   PIN FE_OFN13687_n_143426
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.698 249.792 11.726 ;
      END
   END FE_OFN13687_n_143426

   PIN FE_OFN13692_n_41993
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.33 249.792 57.358 ;
      END
   END FE_OFN13692_n_41993

   PIN FE_OFN14071_n_142964
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.818 0.0 24.846 0.163 ;
      END
   END FE_OFN14071_n_142964

   PIN FE_OFN14164_n_31516
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.698 117.597 43.726 117.76 ;
      END
   END FE_OFN14164_n_31516

   PIN FE_OFN14397_n_140213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.426 249.792 77.454 ;
      END
   END FE_OFN14397_n_140213

   PIN FE_OFN14901_n_140203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 23.41 249.792 23.438 ;
      END
   END FE_OFN14901_n_140203

   PIN FE_OFN15072_n_29125
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.73 117.597 135.758 117.76 ;
      END
   END FE_OFN15072_n_29125

   PIN FE_OFN15106_n_30279
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.634 117.597 139.662 117.76 ;
      END
   END FE_OFN15106_n_30279

   PIN FE_OFN15135_n_30145
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 185.714 117.597 185.742 117.76 ;
      END
   END FE_OFN15135_n_30145

   PIN FE_OFN15329_n_29953
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.954 117.597 131.982 117.76 ;
      END
   END FE_OFN15329_n_29953

   PIN FE_OFN15343_n_30559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.346 117.597 143.374 117.76 ;
      END
   END FE_OFN15343_n_30559

   PIN FE_OFN16079_n_41709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.098 249.792 26.126 ;
      END
   END FE_OFN16079_n_41709

   PIN FE_OFN16087_n_41993
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.026 249.792 55.054 ;
      END
   END FE_OFN16087_n_41993

   PIN FE_OFN16127_n_66979
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 53.426 249.792 53.454 ;
      END
   END FE_OFN16127_n_66979

   PIN FE_OFN16313_b_7_6_9
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.242 249.792 48.27 ;
      END
   END FE_OFN16313_b_7_6_9

   PIN FE_OFN17006_n_58282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.53 117.597 124.558 117.76 ;
      END
   END FE_OFN17006_n_58282

   PIN FE_OFN17423_n_8249
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.018 0.0 228.046 0.163 ;
      END
   END FE_OFN17423_n_8249

   PIN FE_OFN17844_n_81895
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.562 249.792 80.59 ;
      END
   END FE_OFN17844_n_81895

   PIN FE_OFN17850_n_66751
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.018 249.792 84.046 ;
      END
   END FE_OFN17850_n_66751

   PIN FE_OFN17864_n_71795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.322 249.792 30.35 ;
      END
   END FE_OFN17864_n_71795

   PIN FE_OFN17908_n_55576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.65 249.792 49.678 ;
      END
   END FE_OFN17908_n_55576

   PIN FE_OFN18784_n_31306
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.602 117.597 111.63 117.76 ;
      END
   END FE_OFN18784_n_31306

   PIN FE_OFN19276_n_28640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.41 117.597 143.438 117.76 ;
      END
   END FE_OFN19276_n_28640

   PIN FE_OFN2321_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 143.538 117.597 143.566 117.76 ;
      END
   END FE_OFN2321_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_14_

   PIN FE_OFN2322_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 147.378 117.597 147.406 117.76 ;
      END
   END FE_OFN2322_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_13_

   PIN FE_OFN4459_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.322 0.0 142.35 0.163 ;
      END
   END FE_OFN4459_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_12_

   PIN FE_OFN4762_n_137230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.002 0.0 78.03 0.082 ;
      END
   END FE_OFN4762_n_137230

   PIN FE_OFN4815_n_143202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.674 0.0 66.702 0.163 ;
      END
   END FE_OFN4815_n_143202

   PIN FE_OFN6162_delay_mul_ln34_unr7_unr8_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.114 0.0 176.142 0.163 ;
      END
   END FE_OFN6162_delay_mul_ln34_unr7_unr8_stage2_stallmux_z_13_

   PIN FE_OFN6326_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 40.69 249.792 40.718 ;
      END
   END FE_OFN6326_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_7_

   PIN FE_OFN6445_n_64478
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 72.818 249.792 72.846 ;
      END
   END FE_OFN6445_n_64478

   PIN FE_OFN6458_n_59534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.906 249.792 41.934 ;
      END
   END FE_OFN6458_n_59534

   PIN FE_OFN6491_n_41960
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 6.642 249.792 6.67 ;
      END
   END FE_OFN6491_n_41960

   PIN FE_OFN6549_n_41963
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 73.266 249.792 73.294 ;
      END
   END FE_OFN6549_n_41963

   PIN FE_OFN6605_n_140234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.01 249.792 65.038 ;
      END
   END FE_OFN6605_n_140234

   PIN FE_OFN6626_n_41612
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.874 249.792 45.902 ;
      END
   END FE_OFN6626_n_41612

   PIN FE_OFN6749_n_41995
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.65 249.792 33.678 ;
      END
   END FE_OFN6749_n_41995

   PIN FE_OFN6841_n_41015
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.738 249.792 26.766 ;
      END
   END FE_OFN6841_n_41015

   PIN FE_OFN6859_n_143629
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.066 249.792 38.094 ;
      END
   END FE_OFN6859_n_143629

   PIN FE_OFN8170_n_26637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.874 117.597 85.902 117.76 ;
      END
   END FE_OFN8170_n_26637

   PIN FE_OFN8330_n_31307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.362 117.597 181.39 117.76 ;
      END
   END FE_OFN8330_n_31307

   PIN FE_OFN8366_n_31480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.818 117.597 16.846 117.76 ;
      END
   END FE_OFN8366_n_31480

   PIN FE_OFN8464_n_25371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.914 117.597 204.942 117.76 ;
      END
   END FE_OFN8464_n_25371

   PIN FE_OFN8492_n_29557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.082 117.597 132.11 117.76 ;
      END
   END FE_OFN8492_n_29557

   PIN FE_OFN8498_n_28380
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.698 117.597 139.726 117.76 ;
      END
   END FE_OFN8498_n_28380

   PIN FE_OFN8499_n_27857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.274 117.597 124.302 117.76 ;
      END
   END FE_OFN8499_n_27857

   PIN FE_OFN8578_n_29968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.954 249.792 3.982 ;
      END
   END FE_OFN8578_n_29968

   PIN FE_OFN8704_n_31118
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.602 249.792 103.63 ;
      END
   END FE_OFN8704_n_31118

   PIN FE_OFN8719_n_25376
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.274 249.792 92.302 ;
      END
   END FE_OFN8719_n_25376

   PIN FE_OFN9239_delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.666 249.792 103.694 ;
      END
   END FE_OFN9239_delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_

   PIN FE_OFN9472_b_7_8_8
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.994 249.792 27.022 ;
      END
   END FE_OFN9472_b_7_8_8

   PIN FE_OFN9474_b_7_8_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 38.386 249.792 38.414 ;
      END
   END FE_OFN9474_b_7_8_7

   PIN FE_OFN9536_b_7_6_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 61.298 249.792 61.326 ;
      END
   END FE_OFN9536_b_7_6_15

   PIN FE_OFN9540_b_7_6_14
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.698 249.792 99.726 ;
      END
   END FE_OFN9540_b_7_6_14

   PIN FE_OFN9548_b_7_6_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 58.034 249.792 58.062 ;
      END
   END FE_OFN9548_b_7_6_11

   PIN FE_OFN9549_b_7_6_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.778 249.792 57.806 ;
      END
   END FE_OFN9549_b_7_6_10

   PIN FE_OFN9558_b_7_6_6
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 54.834 249.792 54.862 ;
      END
   END FE_OFN9558_b_7_6_6

   PIN FE_OFN9564_b_7_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 88.434 249.792 88.462 ;
      END
   END FE_OFN9564_b_7_6_4

   PIN FE_OFN9577_b_7_6_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.71 49.33 249.792 49.358 ;
      END
   END FE_OFN9577_b_7_6_1

   PIN FE_OFN9879_b_4_8_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.346 0.0 95.374 0.163 ;
      END
   END FE_OFN9879_b_4_8_3

   PIN delay_mul_ln34_unr4_unr2_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.842 0.0 145.87 0.163 ;
      END
   END delay_mul_ln34_unr4_unr2_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr4_unr2_stage2_stallmux_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.778 0.0 65.806 0.163 ;
      END
   END delay_mul_ln34_unr4_unr2_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr4_unr4_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.074 0.0 113.102 0.163 ;
      END
   END delay_mul_ln34_unr4_unr4_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr4_unr6_stage2_stallmux_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 125.426 0.0 125.454 0.163 ;
      END
   END delay_mul_ln34_unr4_unr6_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr4_unr6_stage2_stallmux_z_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.61 0.0 114.638 0.163 ;
      END
   END delay_mul_ln34_unr4_unr6_stage2_stallmux_z_8_

   PIN delay_mul_ln34_unr7_unr0_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 85.234 249.792 85.262 ;
      END
   END delay_mul_ln34_unr7_unr0_stage2_stallmux_q_12_

   PIN delay_mul_ln34_unr7_unr8_stage2_stallmux_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.162 0.0 154.19 0.163 ;
      END
   END delay_mul_ln34_unr7_unr8_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.594 117.597 116.622 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.434 117.597 120.462 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_q_3_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.818 117.597 208.846 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_12_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.498 117.597 120.526 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_4_

   PIN mul_4647_72_n_200
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.082 0.0 4.11 0.163 ;
      END
   END mul_4647_72_n_200

   PIN mul_4647_72_n_224
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.274 0.0 28.302 0.163 ;
      END
   END mul_4647_72_n_224

   PIN mul_4647_72_n_227
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.53 0.0 20.558 0.163 ;
      END
   END mul_4647_72_n_227

   PIN mul_4647_72_n_230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.146 0.0 20.174 0.163 ;
      END
   END mul_4647_72_n_230

   PIN mul_4647_72_n_252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.794 0.0 39.822 0.163 ;
      END
   END mul_4647_72_n_252

   PIN mul_4647_72_n_323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.85 0.0 36.878 0.163 ;
      END
   END mul_4647_72_n_323

   PIN mul_4647_72_n_71
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.978 0.0 13.006 0.163 ;
      END
   END mul_4647_72_n_71

   PIN mul_4649_72_n_77
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.722 0.0 116.75 0.163 ;
      END
   END mul_4649_72_n_77

   PIN mul_4651_72_n_290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.386 0.0 78.414 0.163 ;
      END
   END mul_4651_72_n_290

   PIN mul_4651_72_n_316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.61 0.0 66.638 0.163 ;
      END
   END mul_4651_72_n_316

   PIN mul_4651_72_n_322
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.386 0.0 70.414 0.163 ;
      END
   END mul_4651_72_n_322

   PIN mul_4651_72_n_323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.834 0.0 70.862 0.163 ;
      END
   END mul_4651_72_n_323

   PIN mul_4651_72_n_324
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.282 0.0 71.31 0.163 ;
      END
   END mul_4651_72_n_324

   PIN mul_4664_72_n_213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.114 0.0 32.142 0.163 ;
      END
   END mul_4664_72_n_213

   PIN mul_4664_72_n_214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.178 0.0 32.206 0.163 ;
      END
   END mul_4664_72_n_214

   PIN mul_4664_72_n_285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.402 0.0 28.43 0.163 ;
      END
   END mul_4664_72_n_285

   PIN mul_4664_72_n_55
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 0.0 25.614 0.163 ;
      END
   END mul_4664_72_n_55

   PIN mul_4664_72_n_71
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.522 0.0 25.55 0.163 ;
      END
   END mul_4664_72_n_71

   PIN mul_4664_72_n_773
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.05 0.0 32.078 0.163 ;
      END
   END mul_4664_72_n_773

   PIN mul_4698_72_n_117
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.13 249.792 38.158 ;
      END
   END mul_4698_72_n_117

   PIN mul_4700_72_n_53
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 4.146 249.792 4.174 ;
      END
   END mul_4700_72_n_53

   PIN mul_4700_72_n_69
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 4.21 249.792 4.238 ;
      END
   END mul_4700_72_n_69

   PIN n_100733
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.234 117.597 197.262 117.76 ;
      END
   END n_100733

   PIN n_100744
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 189.682 117.597 189.71 117.76 ;
      END
   END n_100744

   PIN n_102607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 61.17 249.792 61.198 ;
      END
   END n_102607

   PIN n_102890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.282 0.0 151.31 0.163 ;
      END
   END n_102890

   PIN n_103077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.298 117.597 197.326 117.76 ;
      END
   END n_103077

   PIN n_103482
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 212.658 117.597 212.686 117.76 ;
      END
   END n_103482

   PIN n_105239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.722 117.597 212.75 117.76 ;
      END
   END n_105239

   PIN n_106473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 189.49 117.597 189.518 117.76 ;
      END
   END n_106473

   PIN n_107990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.266 0.0 41.294 0.163 ;
      END
   END n_107990

   PIN n_108077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.706 117.597 182.734 117.76 ;
      END
   END n_108077

   PIN n_108091
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.138 117.597 201.166 117.76 ;
      END
   END n_108091

   PIN n_108970
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.626 0.0 40.654 0.163 ;
      END
   END n_108970

   PIN n_109766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.634 117.597 203.662 117.76 ;
      END
   END n_109766

   PIN n_110534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 183.986 117.597 184.014 117.76 ;
      END
   END n_110534

   PIN n_110678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.074 249.792 65.102 ;
      END
   END n_110678

   PIN n_110705
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.658 117.597 180.686 117.76 ;
      END
   END n_110705

   PIN n_11212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.962 0.0 14.99 0.163 ;
      END
   END n_11212

   PIN n_11214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.714 249.792 49.742 ;
      END
   END n_11214

   PIN n_114514
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.306 0.0 32.334 0.163 ;
      END
   END n_114514

   PIN n_115085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.186 0.0 35.214 0.163 ;
      END
   END n_115085

   PIN n_115534
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.258 117.597 54.286 117.76 ;
      END
   END n_115534

   PIN n_115535
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.818 117.597 48.846 117.76 ;
      END
   END n_115535

   PIN n_115594
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.786 0.0 20.814 0.163 ;
      END
   END n_115594

   PIN n_115658
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 51.25 0.0 51.278 0.163 ;
      END
   END n_115658

   PIN n_116050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.018 0.0 44.046 0.163 ;
      END
   END n_116050

   PIN n_116051
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.018 0.0 44.046 0.163 ;
      END
   END n_116051

   PIN n_116348
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.346 0.0 47.374 0.163 ;
      END
   END n_116348

   PIN n_116462
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.698 0.0 3.726 0.163 ;
      END
   END n_116462

   PIN n_116511
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.026 0.0 55.054 0.163 ;
      END
   END n_116511

   PIN n_116767
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.178 0.0 32.206 0.163 ;
      END
   END n_116767

   PIN n_116839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.842 0.0 41.87 0.163 ;
      END
   END n_116839

   PIN n_118700
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.442 0.0 3.47 0.163 ;
      END
   END n_118700

   PIN n_118762
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.258 0.0 22.286 0.163 ;
      END
   END n_118762

   PIN n_118773
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.042 0.0 5.07 0.163 ;
      END
   END n_118773

   PIN n_118968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.69 0.0 16.718 0.163 ;
      END
   END n_118968

   PIN n_118969
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.786 0.0 12.814 0.163 ;
      END
   END n_118969

   PIN n_118970
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.042 0.0 13.07 0.163 ;
      END
   END n_118970

   PIN n_119000
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.89 0.0 43.918 0.163 ;
      END
   END n_119000

   PIN n_119073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.034 117.597 10.062 117.76 ;
      END
   END n_119073

   PIN n_119481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.546 0.0 18.574 0.163 ;
      END
   END n_119481

   PIN n_119509
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.538 0.0 47.566 0.163 ;
      END
   END n_119509

   PIN n_120297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.802 0.0 10.83 0.163 ;
      END
   END n_120297

   PIN n_120453
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.242 0.0 32.27 0.163 ;
      END
   END n_120453

   PIN n_120804
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.37 0.0 48.398 0.163 ;
      END
   END n_120804

   PIN n_120838
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.506 0.0 3.534 0.163 ;
      END
   END n_120838

   PIN n_120840
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.994 0.0 19.022 0.163 ;
      END
   END n_120840

   PIN n_121307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.194 0.0 78.222 0.163 ;
      END
   END n_121307

   PIN n_121492
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.338 0.0 28.366 0.163 ;
      END
   END n_121492

   PIN n_121670
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.226 0.0 74.254 0.163 ;
      END
   END n_121670

   PIN n_121988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.434 0.0 24.462 0.163 ;
      END
   END n_121988

   PIN n_122043
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.442 117.597 3.47 117.76 ;
      END
   END n_122043

   PIN n_122081
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.626 0.0 24.654 0.163 ;
      END
   END n_122081

   PIN n_122221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.786 0.0 4.814 0.163 ;
      END
   END n_122221

   PIN n_122483
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.666 0.163 7.694 ;
      END
   END n_122483

   PIN n_122484
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.282 0.163 55.31 ;
      END
   END n_122484

   PIN n_122506
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.306 117.597 8.334 117.76 ;
      END
   END n_122506

   PIN n_122507
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.786 117.597 4.814 117.76 ;
      END
   END n_122507

   PIN n_123326
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.138 0.0 9.166 0.163 ;
      END
   END n_123326

   PIN n_124275
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.362 0.0 5.39 0.163 ;
      END
   END n_124275

   PIN n_124317
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.466 0.0 20.494 0.163 ;
      END
   END n_124317

   PIN n_124544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.81 117.597 37.838 117.76 ;
      END
   END n_124544

   PIN n_124640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.954 117.597 51.982 117.76 ;
      END
   END n_124640

   PIN n_124871
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.594 0.0 20.622 0.163 ;
      END
   END n_124871

   PIN n_126137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.794 117.597 39.822 117.76 ;
      END
   END n_126137

   PIN n_127194
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.85 0.0 12.878 0.163 ;
      END
   END n_127194

   PIN n_127226
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.954 117.597 35.982 117.76 ;
      END
   END n_127226

   PIN n_127725
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.57 0.0 3.598 0.163 ;
      END
   END n_127725

   PIN n_127726
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.554 0.0 5.582 0.163 ;
      END
   END n_127726

   PIN n_128154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.658 0.0 28.686 0.163 ;
      END
   END n_128154

   PIN n_128155
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.658 0.0 20.686 0.163 ;
      END
   END n_128155

   PIN n_128174
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.306 0.0 24.334 0.163 ;
      END
   END n_128174

   PIN n_128290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.914 0.0 12.942 0.163 ;
      END
   END n_128290

   PIN n_128294
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.714 0.0 9.742 0.163 ;
      END
   END n_128294

   PIN n_129242
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.106 117.597 21.134 117.76 ;
      END
   END n_129242

   PIN n_129244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.762 117.597 27.79 117.76 ;
      END
   END n_129244

   PIN n_129371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.226 0.163 114.254 ;
      END
   END n_129371

   PIN n_129623
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.394 0.0 9.422 0.163 ;
      END
   END n_129623

   PIN n_129649
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.762 0.163 3.79 ;
      END
   END n_129649

   PIN n_129721
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.266 0.0 9.294 0.163 ;
      END
   END n_129721

   PIN n_130485
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.69 117.597 24.718 117.76 ;
      END
   END n_130485

   PIN n_131556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.562 117.597 32.59 117.76 ;
      END
   END n_131556

   PIN n_133552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.978 0.0 37.006 0.163 ;
      END
   END n_133552

   PIN n_134508
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.162 0.0 18.19 0.163 ;
      END
   END n_134508

   PIN n_135085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.754 0.0 16.782 0.163 ;
      END
   END n_135085

   PIN n_137235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 38.322 249.792 38.35 ;
      END
   END n_137235

   PIN n_137837
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.37 0.0 88.398 0.163 ;
      END
   END n_137837

   PIN n_143371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.09 249.792 15.118 ;
      END
   END n_143371

   PIN n_143818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.53 0.0 12.558 0.163 ;
      END
   END n_143818

   PIN n_24537
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 194.802 0.0 194.83 0.163 ;
      END
   END n_24537

   PIN n_24538
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 193.33 0.0 193.358 0.163 ;
      END
   END n_24538

   PIN n_25880
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 171.186 0.0 171.214 0.163 ;
      END
   END n_25880

   PIN n_25882
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.354 0.0 170.382 0.163 ;
      END
   END n_25882

   PIN n_26382
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.314 117.597 147.342 117.76 ;
      END
   END n_26382

   PIN n_26770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.498 117.597 144.526 117.76 ;
      END
   END n_26770

   PIN n_26771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 147.314 117.597 147.342 117.76 ;
      END
   END n_26771

   PIN n_26989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 4.594 249.792 4.622 ;
      END
   END n_26989

   PIN n_27355
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.986 117.597 104.014 117.76 ;
      END
   END n_27355

   PIN n_28369
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.89 117.597 131.918 117.76 ;
      END
   END n_28369

   PIN n_2842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.61 0.0 10.638 0.163 ;
      END
   END n_2842

   PIN n_28483
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.754 117.597 208.782 117.76 ;
      END
   END n_28483

   PIN n_28878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 178.098 117.597 178.126 117.76 ;
      END
   END n_28878

   PIN n_29113
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.858 249.792 103.886 ;
      END
   END n_29113

   PIN n_2937
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.586 0.0 121.614 0.163 ;
      END
   END n_2937

   PIN n_29558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.018 117.597 132.046 117.76 ;
      END
   END n_29558

   PIN n_32569
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.282 0.0 47.31 0.163 ;
      END
   END n_32569

   PIN n_32599
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.378 0.0 67.406 0.163 ;
      END
   END n_32599

   PIN n_32677
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.954 0.0 75.982 0.163 ;
      END
   END n_32677

   PIN n_32709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.098 0.0 50.126 0.163 ;
      END
   END n_32709

   PIN n_32886
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.73 0.0 39.758 0.163 ;
      END
   END n_32886

   PIN n_33168
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 19.25 249.792 19.278 ;
      END
   END n_33168

   PIN n_33209
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.09 0.0 55.118 0.163 ;
      END
   END n_33209

   PIN n_33371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.626 249.792 40.654 ;
      END
   END n_33371

   PIN n_34045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.498 0.0 24.526 0.163 ;
      END
   END n_34045

   PIN n_34363
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.65 0.0 81.678 0.163 ;
      END
   END n_34363

   PIN n_34386
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.626 0.0 112.654 0.163 ;
      END
   END n_34386

   PIN n_34739
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.578 249.792 22.606 ;
      END
   END n_34739

   PIN n_35423
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.586 0.0 81.614 0.163 ;
      END
   END n_35423

   PIN n_36289
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.154 0.0 71.182 0.163 ;
      END
   END n_36289

   PIN n_36486
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.322 0.0 78.35 0.163 ;
      END
   END n_36486

   PIN n_36699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.098 0.0 58.126 0.163 ;
      END
   END n_36699

   PIN n_36728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.962 0.0 70.99 0.163 ;
      END
   END n_36728

   PIN n_36741
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.986 249.792 8.014 ;
      END
   END n_36741

   PIN n_36776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 53.874 249.792 53.902 ;
      END
   END n_36776

   PIN n_36951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.57 0.0 43.598 0.163 ;
      END
   END n_36951

   PIN n_37371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.794 0.0 39.822 0.163 ;
      END
   END n_37371

   PIN n_37496
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.634 0.0 75.662 0.163 ;
      END
   END n_37496

   PIN n_37823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.162 0.0 74.19 0.163 ;
      END
   END n_37823

   PIN n_38020
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.626 0.0 64.654 0.163 ;
      END
   END n_38020

   PIN n_38377
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.042 0.0 37.07 0.163 ;
      END
   END n_38377

   PIN n_39631
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.602 0.0 39.63 0.163 ;
      END
   END n_39631

   PIN n_40828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.81 249.792 37.838 ;
      END
   END n_40828

   PIN n_40903
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.706 0.0 70.734 0.163 ;
      END
   END n_40903

   PIN n_43135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.842 117.597 241.87 117.76 ;
      END
   END n_43135

   PIN n_43460
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.042 249.792 77.07 ;
      END
   END n_43460

   PIN n_43886
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.962 249.792 30.99 ;
      END
   END n_43886

   PIN n_43887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.578 249.792 30.606 ;
      END
   END n_43887

   PIN n_43927
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.49 249.792 77.518 ;
      END
   END n_43927

   PIN n_43959
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.314 249.792 11.342 ;
      END
   END n_43959

   PIN n_44225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.17 249.792 77.198 ;
      END
   END n_44225

   PIN n_44595
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.698 117.597 235.726 117.76 ;
      END
   END n_44595

   PIN n_44641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.642 249.792 22.67 ;
      END
   END n_44641

   PIN n_44714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.394 249.792 57.422 ;
      END
   END n_44714

   PIN n_44715
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.714 249.792 57.742 ;
      END
   END n_44715

   PIN n_44776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.874 249.792 37.902 ;
      END
   END n_44776

   PIN n_44777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.258 249.792 38.286 ;
      END
   END n_44777

   PIN n_45142
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 34.226 249.792 34.254 ;
      END
   END n_45142

   PIN n_45217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.626 249.792 80.654 ;
      END
   END n_45217

   PIN n_45222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.954 0.0 131.982 0.163 ;
      END
   END n_45222

   PIN n_45299
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 178.034 0.0 178.062 0.163 ;
      END
   END n_45299

   PIN n_45510
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.53 0.0 116.558 0.163 ;
      END
   END n_45510

   PIN n_45631
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.01 0.0 81.038 0.163 ;
      END
   END n_45631

   PIN n_45632
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.074 0.0 81.102 0.163 ;
      END
   END n_45632

   PIN n_45699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 34.29 249.792 34.318 ;
      END
   END n_45699

   PIN n_45883
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.554 249.792 77.582 ;
      END
   END n_45883

   PIN n_46067
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.018 0.0 132.046 0.163 ;
      END
   END n_46067

   PIN n_46081
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.282 249.792 55.31 ;
      END
   END n_46081

   PIN n_46203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 178.098 0.0 178.126 0.163 ;
      END
   END n_46203

   PIN n_46332
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.562 249.792 48.59 ;
      END
   END n_46332

   PIN n_46335
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 249.01 0.0 249.038 0.163 ;
      END
   END n_46335

   PIN n_46361
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.842 249.792 41.87 ;
      END
   END n_46361

   PIN n_46369
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 85.362 249.792 85.39 ;
      END
   END n_46369

   PIN n_46370
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 85.618 249.792 85.646 ;
      END
   END n_46370

   PIN n_46467
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 80.626 249.792 80.654 ;
      END
   END n_46467

   PIN n_46468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 99.762 249.792 99.79 ;
      END
   END n_46468

   PIN n_46540
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 53.234 249.792 53.262 ;
      END
   END n_46540

   PIN n_46576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.618 0.0 117.646 0.163 ;
      END
   END n_46576

   PIN n_46582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.522 249.792 65.55 ;
      END
   END n_46582

   PIN n_46583
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.178 0.0 224.206 0.163 ;
      END
   END n_46583

   PIN n_46659
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.378 249.792 11.406 ;
      END
   END n_46659

   PIN n_46661
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.354 0.0 114.382 0.163 ;
      END
   END n_46661

   PIN n_46668
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.522 249.792 49.55 ;
      END
   END n_46668

   PIN n_46669
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.33 249.792 49.358 ;
      END
   END n_46669

   PIN n_46676
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 58.354 249.792 58.382 ;
      END
   END n_46676

   PIN n_46872
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.458 249.792 57.486 ;
      END
   END n_46872

   PIN n_46916
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.898 0.0 94.926 0.163 ;
      END
   END n_46916

   PIN n_46917
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.994 0.0 83.022 0.163 ;
      END
   END n_46917

   PIN n_47149
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.778 249.792 49.806 ;
      END
   END n_47149

   PIN n_47248
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 88.498 249.792 88.526 ;
      END
   END n_47248

   PIN n_47260
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.698 0.0 139.726 0.163 ;
      END
   END n_47260

   PIN n_47323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.874 0.0 181.902 0.163 ;
      END
   END n_47323

   PIN n_47423
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 85.426 249.792 85.454 ;
      END
   END n_47423

   PIN n_47856
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.506 0.0 51.534 0.163 ;
      END
   END n_47856

   PIN n_47857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.122 0.0 51.15 0.163 ;
      END
   END n_47857

   PIN n_49211
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.858 0.0 31.886 0.163 ;
      END
   END n_49211

   PIN n_49947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.386 249.792 30.414 ;
      END
   END n_49947

   PIN n_50245
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 88.242 249.792 88.27 ;
      END
   END n_50245

   PIN n_50316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 236.786 117.597 236.814 117.76 ;
      END
   END n_50316

   PIN n_50589
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.298 249.792 77.326 ;
      END
   END n_50589

   PIN n_50941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.858 249.792 47.886 ;
      END
   END n_50941

   PIN n_51049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.906 0.0 129.934 0.163 ;
      END
   END n_51049

   PIN n_51080
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.81 0.0 181.838 0.163 ;
      END
   END n_51080

   PIN n_51152
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.298 0.0 109.326 0.163 ;
      END
   END n_51152

   PIN n_51247
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 54.962 249.792 54.99 ;
      END
   END n_51247

   PIN n_52208
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.194 249.792 38.222 ;
      END
   END n_52208

   PIN n_52412
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.138 249.792 65.166 ;
      END
   END n_52412

   PIN n_52666
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 61.17 249.792 61.198 ;
      END
   END n_52666

   PIN n_52803
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 85.49 249.792 85.518 ;
      END
   END n_52803

   PIN n_52852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.634 117.597 235.662 117.76 ;
      END
   END n_52852

   PIN n_53092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.634 0.0 139.662 0.163 ;
      END
   END n_53092

   PIN n_53255
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 88.306 249.792 88.334 ;
      END
   END n_53255

   PIN n_53257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 42.034 249.792 42.062 ;
      END
   END n_53257

   PIN n_53297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.45 249.792 70.478 ;
      END
   END n_53297

   PIN n_53524
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.578 249.792 38.606 ;
      END
   END n_53524

   PIN n_53555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.826 249.792 99.854 ;
      END
   END n_53555

   PIN n_53566
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.834 117.597 246.862 117.76 ;
      END
   END n_53566

   PIN n_53983
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.738 0.0 82.766 0.163 ;
      END
   END n_53983

   PIN n_53996
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 53.49 249.792 53.518 ;
      END
   END n_53996

   PIN n_54311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.154 0.0 55.182 0.163 ;
      END
   END n_54311

   PIN n_54338
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.362 249.792 77.39 ;
      END
   END n_54338

   PIN n_54688
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.45 249.792 30.478 ;
      END
   END n_54688

   PIN n_54944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.794 117.597 135.822 117.76 ;
      END
   END n_54944

   PIN n_54954
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.314 117.597 115.342 117.76 ;
      END
   END n_54954

   PIN n_54986
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 236.658 117.597 236.686 117.76 ;
      END
   END n_54986

   PIN n_55042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.018 249.792 92.046 ;
      END
   END n_55042

   PIN n_55157
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.386 117.597 158.414 117.76 ;
      END
   END n_55157

   PIN n_55513
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 34.354 249.792 34.382 ;
      END
   END n_55513

   PIN n_5555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 9.01 249.792 9.038 ;
      END
   END n_5555

   PIN n_55597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.266 249.792 41.294 ;
      END
   END n_55597

   PIN n_55598
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.514 249.792 30.542 ;
      END
   END n_55598

   PIN n_55674
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 174.194 0.0 174.222 0.163 ;
      END
   END n_55674

   PIN n_55702
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.93 0.0 58.958 0.163 ;
      END
   END n_55702

   PIN n_55723
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.57 0.0 139.598 0.163 ;
      END
   END n_55723

   PIN n_55740
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.93 0.0 154.958 0.163 ;
      END
   END n_55740

   PIN n_55766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.586 249.792 33.614 ;
      END
   END n_55766

   PIN n_56659
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.202 249.792 65.23 ;
      END
   END n_56659

   PIN n_56808
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.082 249.792 92.11 ;
      END
   END n_56808

   PIN n_56899
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 85.298 249.792 85.326 ;
      END
   END n_56899

   PIN n_57040
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.762 0.0 83.79 0.163 ;
      END
   END n_57040

   PIN n_57135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.826 0.163 3.854 ;
      END
   END n_57135

   PIN n_57460
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.714 0.0 137.742 0.163 ;
      END
   END n_57460

   PIN n_57673
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 183.346 0.0 183.374 0.163 ;
      END
   END n_57673

   PIN n_57704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.642 249.792 38.67 ;
      END
   END n_57704

   PIN n_57712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.442 0.0 163.47 0.163 ;
      END
   END n_57712

   PIN n_57713
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.738 0.0 162.766 0.163 ;
      END
   END n_57713

   PIN n_57714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.122 0.0 163.15 0.163 ;
      END
   END n_57714

   PIN n_57823
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 58.226 249.792 58.254 ;
      END
   END n_57823

   PIN n_57902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.69 117.597 112.718 117.76 ;
      END
   END n_57902

   PIN n_57982
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 158.898 117.597 158.926 117.76 ;
      END
   END n_57982

   PIN n_58071
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.938 249.792 45.966 ;
      END
   END n_58071

   PIN n_58207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.706 249.792 38.734 ;
      END
   END n_58207

   PIN n_58229
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.794 117.597 231.822 117.76 ;
      END
   END n_58229

   PIN n_58234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 178.162 117.597 178.19 117.76 ;
      END
   END n_58234

   PIN n_58257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.098 117.597 162.126 117.76 ;
      END
   END n_58257

   PIN n_58264
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.85 117.597 132.878 117.76 ;
      END
   END n_58264

   PIN n_58283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.21 117.597 124.238 117.76 ;
      END
   END n_58283

   PIN n_58292
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.474 0.0 143.502 0.163 ;
      END
   END n_58292

   PIN n_58507
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 46.002 249.792 46.03 ;
      END
   END n_58507

   PIN n_59057
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.946 117.597 152.974 117.76 ;
      END
   END n_59057

   PIN n_59287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.77 117.597 158.798 117.76 ;
      END
   END n_59287

   PIN n_59495
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 155.058 0.0 155.086 0.163 ;
      END
   END n_59495

   PIN n_59615
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.866 249.792 106.894 ;
      END
   END n_59615

   PIN n_59894
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.634 0.0 3.662 0.163 ;
      END
   END n_59894

   PIN n_60087
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 236.402 117.597 236.43 117.76 ;
      END
   END n_60087

   PIN n_60088
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 135.858 117.597 135.886 117.76 ;
      END
   END n_60088

   PIN n_60104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.666 249.792 47.694 ;
      END
   END n_60104

   PIN n_60139
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.146 249.792 92.174 ;
      END
   END n_60139

   PIN n_60261
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 95.986 249.792 96.014 ;
      END
   END n_60261

   PIN n_60264
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.026 117.597 159.054 117.76 ;
      END
   END n_60264

   PIN n_60317
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.002 117.597 126.03 117.76 ;
      END
   END n_60317

   PIN n_60318
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.066 117.597 126.094 117.76 ;
      END
   END n_60318

   PIN n_60377
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 72.69 249.792 72.718 ;
      END
   END n_60377

   PIN n_60444
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.73 249.792 103.758 ;
      END
   END n_60444

   PIN n_60543
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.498 249.792 48.526 ;
      END
   END n_60543

   PIN n_60569
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 178.162 0.0 178.19 0.163 ;
      END
   END n_60569

   PIN n_60575
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.378 0.0 163.406 0.163 ;
      END
   END n_60575

   PIN n_60581
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.754 0.0 176.782 0.163 ;
      END
   END n_60581

   PIN n_60661
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.138 117.597 113.166 117.76 ;
      END
   END n_60661

   PIN n_60763
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 31.474 249.792 31.502 ;
      END
   END n_60763

   PIN n_60770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.138 117.597 137.166 117.76 ;
      END
   END n_60770

   PIN n_61110
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.938 117.597 85.966 117.76 ;
      END
   END n_61110

   PIN n_61151
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.306 0.0 112.334 0.163 ;
      END
   END n_61151

   PIN n_61597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.842 249.792 57.87 ;
      END
   END n_61597

   PIN n_61600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 53.298 249.792 53.326 ;
      END
   END n_61600

   PIN n_61622
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.834 0.0 158.862 0.163 ;
      END
   END n_61622

   PIN n_61766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.714 0.0 89.742 0.163 ;
      END
   END n_61766

   PIN n_61876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.754 117.597 160.782 117.76 ;
      END
   END n_61876

   PIN n_61877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.61 117.597 162.638 117.76 ;
      END
   END n_61877

   PIN n_61881
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.866 117.597 154.894 117.76 ;
      END
   END n_61881

   PIN n_61896
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.522 117.597 129.55 117.76 ;
      END
   END n_61896

   PIN n_62357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.186 117.597 91.214 117.76 ;
      END
   END n_62357

   PIN n_62360
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.474 249.792 15.502 ;
      END
   END n_62360

   PIN n_62401
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.394 0.0 105.422 0.163 ;
      END
   END n_62401

   PIN n_62504
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.138 249.792 41.166 ;
      END
   END n_62504

   PIN n_62647
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.146 117.597 164.174 117.76 ;
      END
   END n_62647

   PIN n_62807
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.338 117.597 68.366 117.76 ;
      END
   END n_62807

   PIN n_62808
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.474 117.597 71.502 117.76 ;
      END
   END n_62808

   PIN n_62998
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.522 117.597 97.55 117.76 ;
      END
   END n_62998

   PIN n_63006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.778 249.792 33.806 ;
      END
   END n_63006

   PIN n_63048
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 73.01 249.792 73.038 ;
      END
   END n_63048

   PIN n_63049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 73.074 249.792 73.102 ;
      END
   END n_63049

   PIN n_63050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.442 0.0 155.47 0.163 ;
      END
   END n_63050

   PIN n_63051
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.506 0.0 155.534 0.163 ;
      END
   END n_63051

   PIN n_63137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.962 249.792 14.99 ;
      END
   END n_63137

   PIN n_63203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.074 249.792 33.102 ;
      END
   END n_63203

   PIN n_63244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.674 117.597 162.702 117.76 ;
      END
   END n_63244

   PIN n_63246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.858 117.597 135.886 117.76 ;
      END
   END n_63246

   PIN n_63253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 248.498 117.597 248.526 117.76 ;
      END
   END n_63253

   PIN n_63258
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.37 117.597 216.398 117.76 ;
      END
   END n_63258

   PIN n_63272
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.914 0.0 204.942 0.163 ;
      END
   END n_63272

   PIN n_63359
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 185.138 0.0 185.166 0.163 ;
      END
   END n_63359

   PIN n_63530
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 155.058 117.597 155.086 117.76 ;
      END
   END n_63530

   PIN n_63531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 153.074 117.597 153.102 117.76 ;
      END
   END n_63531

   PIN n_63563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.138 117.597 89.166 117.76 ;
      END
   END n_63563

   PIN n_6357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.458 0.0 121.486 0.163 ;
      END
   END n_6357

   PIN n_63724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.538 249.792 15.566 ;
      END
   END n_63724

   PIN n_64400
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.842 249.792 49.87 ;
      END
   END n_64400

   PIN n_64412
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.994 0.0 155.022 0.163 ;
      END
   END n_64412

   PIN n_64413
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.866 0.0 154.894 0.163 ;
      END
   END n_64413

   PIN n_64467
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 99.826 117.597 99.854 117.76 ;
      END
   END n_64467

   PIN n_64527
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 72.946 249.792 72.974 ;
      END
   END n_64527

   PIN n_64551
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.154 117.597 151.182 117.76 ;
      END
   END n_64551

   PIN n_64555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.946 117.597 144.974 117.76 ;
      END
   END n_64555

   PIN n_64556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.762 117.597 147.79 117.76 ;
      END
   END n_64556

   PIN n_64558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.882 117.597 128.91 117.76 ;
      END
   END n_64558

   PIN n_64834
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.538 0.0 143.566 0.163 ;
      END
   END n_64834

   PIN n_64921
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.714 249.792 33.742 ;
      END
   END n_64921

   PIN n_64944
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 72.882 249.792 72.91 ;
      END
   END n_64944

   PIN n_64988
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.57 0.0 91.598 0.163 ;
      END
   END n_64988

   PIN n_65021
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.346 117.597 159.374 117.76 ;
      END
   END n_65021

   PIN n_65147
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.01 117.597 153.038 117.76 ;
      END
   END n_65147

   PIN n_65154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.154 249.792 15.182 ;
      END
   END n_65154

   PIN n_65353
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.922 117.597 143.95 117.76 ;
      END
   END n_65353

   PIN n_65402
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 185.714 0.0 185.742 0.163 ;
      END
   END n_65402

   PIN n_65488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 68.658 249.792 68.686 ;
      END
   END n_65488

   PIN n_65500
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.93 117.597 154.958 117.76 ;
      END
   END n_65500

   PIN n_65528
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.978 0.0 205.006 0.163 ;
      END
   END n_65528

   PIN n_65632
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.25 117.597 155.278 117.76 ;
      END
   END n_65632

   PIN n_65654
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.282 117.597 159.31 117.76 ;
      END
   END n_65654

   PIN n_65680
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.082 0.0 148.11 0.163 ;
      END
   END n_65680

   PIN n_65751
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.33 117.597 153.358 117.76 ;
      END
   END n_65751

   PIN n_65798
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.218 117.597 95.246 117.76 ;
      END
   END n_65798

   PIN n_65952
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.874 0.0 85.902 0.163 ;
      END
   END n_65952

   PIN n_65974
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.762 249.792 11.79 ;
      END
   END n_65974

   PIN n_66586
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.706 249.792 22.734 ;
      END
   END n_66586

   PIN n_66611
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.058 0.0 155.086 0.163 ;
      END
   END n_66611

   PIN n_66722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.882 117.597 224.91 117.76 ;
      END
   END n_66722

   PIN n_66841
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.242 249.792 80.27 ;
      END
   END n_66841

   PIN n_67151
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.186 117.597 155.214 117.76 ;
      END
   END n_67151

   PIN n_67191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.818 117.597 144.846 117.76 ;
      END
   END n_67191

   PIN n_71276
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 31.41 249.792 31.438 ;
      END
   END n_71276

   PIN n_71277
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 31.026 249.792 31.054 ;
      END
   END n_71277

   PIN n_71278
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 31.282 249.792 31.31 ;
      END
   END n_71278

   PIN n_71434
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.066 249.792 30.094 ;
      END
   END n_71434

   PIN n_71435
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.802 249.792 26.83 ;
      END
   END n_71435

   PIN n_71444
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.482 0.0 90.51 0.163 ;
      END
   END n_71444

   PIN n_71763
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 34.418 249.792 34.446 ;
      END
   END n_71763

   PIN n_71770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.306 249.792 80.334 ;
      END
   END n_71770

   PIN n_72006
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.09 117.597 151.118 117.76 ;
      END
   END n_72006

   PIN n_72275
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 68.722 249.792 68.75 ;
      END
   END n_72275

   PIN n_77145
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.122 117.597 155.15 117.76 ;
      END
   END n_77145

   PIN n_77670
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 8.05 249.792 8.078 ;
      END
   END n_77670

   PIN n_77995
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.362 117.597 197.39 117.76 ;
      END
   END n_77995

   PIN n_78280
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.818 249.792 80.846 ;
      END
   END n_78280

   PIN n_78473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.594 117.597 140.622 117.76 ;
      END
   END n_78473

   PIN n_8031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.738 0.0 10.766 0.163 ;
      END
   END n_8031

   PIN n_82565
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.69 249.792 80.718 ;
      END
   END n_82565

   PIN n_83303
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.858 117.597 231.886 117.76 ;
      END
   END n_83303

   PIN n_8403
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 97.458 0.0 97.486 0.163 ;
      END
   END n_8403

   PIN n_84678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.754 249.792 80.782 ;
      END
   END n_84678

   PIN n_85584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.154 0.0 151.182 0.163 ;
      END
   END n_85584

   PIN n_88925
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 96.114 249.792 96.142 ;
      END
   END n_88925

   PIN n_91246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 190.962 117.597 190.99 117.76 ;
      END
   END n_91246

   PIN n_91249
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 247.218 117.597 247.246 117.76 ;
      END
   END n_91249

   PIN n_91279
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.922 117.597 231.95 117.76 ;
      END
   END n_91279

   PIN n_91722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.77 249.792 38.798 ;
      END
   END n_91722

   PIN n_91724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.978 117.597 109.006 117.76 ;
      END
   END n_91724

   PIN n_92857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 23.474 249.792 23.502 ;
      END
   END n_92857

   PIN n_94960
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 96.178 249.792 96.206 ;
      END
   END n_94960

   PIN n_96293
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.57 117.597 139.598 117.76 ;
      END
   END n_96293

   PIN n_97165
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.018 117.597 228.046 117.76 ;
      END
   END n_97165

   PIN n_97291
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.194 0.0 110.222 0.163 ;
      END
   END n_97291

   PIN FE_OFN10008_b_4_4_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.65 0.0 41.678 0.163 ;
      END
   END FE_OFN10008_b_4_4_11

   PIN FE_OFN10010_b_4_4_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 41.97 0.0 41.998 0.163 ;
      END
   END FE_OFN10010_b_4_4_10

   PIN FE_OFN10012_b_4_4_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.434 0.0 48.462 0.163 ;
      END
   END FE_OFN10012_b_4_4_9

   PIN FE_OFN10014_b_4_4_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.834 0.0 14.862 0.163 ;
      END
   END FE_OFN10014_b_4_4_8

   PIN FE_OFN10015_b_4_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.866 0.0 58.894 0.163 ;
      END
   END FE_OFN10015_b_4_4_7

   PIN FE_OFN10022_b_4_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.89 0.0 35.918 0.163 ;
      END
   END FE_OFN10022_b_4_4_5

   PIN FE_OFN10023_b_4_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.362 0.0 37.39 0.163 ;
      END
   END FE_OFN10023_b_4_4_5

   PIN FE_OFN10027_b_4_4_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.986 0.0 32.014 0.163 ;
      END
   END FE_OFN10027_b_4_4_3

   PIN FE_OFN10031_b_4_4_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.602 0.0 47.63 0.163 ;
      END
   END FE_OFN10031_b_4_4_2

   PIN FE_OFN10037_b_4_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.978 0.0 21.006 0.163 ;
      END
   END FE_OFN10037_b_4_4_0

   PIN FE_OFN10082_b_4_2_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.858 0.0 39.886 0.163 ;
      END
   END FE_OFN10082_b_4_2_12

   PIN FE_OFN10084_b_4_2_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.498 0.0 56.526 0.163 ;
      END
   END FE_OFN10084_b_4_2_11

   PIN FE_OFN10086_b_4_2_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.866 0.0 58.894 0.163 ;
      END
   END FE_OFN10086_b_4_2_10

   PIN FE_OFN10088_b_4_2_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.666 0.0 39.694 0.163 ;
      END
   END FE_OFN10088_b_4_2_9

   PIN FE_OFN10090_b_4_2_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.994 0.0 35.022 0.163 ;
      END
   END FE_OFN10090_b_4_2_8

   PIN FE_OFN10093_b_4_2_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.578 0.0 30.606 0.163 ;
      END
   END FE_OFN10093_b_4_2_7

   PIN FE_OFN10098_b_4_2_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.466 0.0 28.494 0.082 ;
      END
   END FE_OFN10098_b_4_2_5

   PIN FE_OFN10100_b_4_2_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.69 0.0 24.718 0.082 ;
      END
   END FE_OFN10100_b_4_2_4

   PIN FE_OFN10102_b_4_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.274 0.0 60.302 0.082 ;
      END
   END FE_OFN10102_b_4_2_3

   PIN FE_OFN10104_b_4_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.754 0.0 24.782 0.163 ;
      END
   END FE_OFN10104_b_4_2_2

   PIN FE_OFN10105_b_4_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.098 0.0 90.126 0.163 ;
      END
   END FE_OFN10105_b_4_2_2

   PIN FE_OFN10106_b_4_2_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.466 0.0 60.494 0.163 ;
      END
   END FE_OFN10106_b_4_2_1

   PIN FE_OFN10110_b_4_2_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.226 0.0 58.254 0.082 ;
      END
   END FE_OFN10110_b_4_2_0

   PIN FE_OFN11414_n_140210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 62.898 249.792 62.926 ;
      END
   END FE_OFN11414_n_140210

   PIN FE_OFN11419_n_140210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.71 15.346 249.792 15.374 ;
      END
   END FE_OFN11419_n_140210

   PIN FE_OFN11481_n_140205
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.994 249.792 19.022 ;
      END
   END FE_OFN11481_n_140205

   PIN FE_OFN11522_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.434 249.792 48.462 ;
      END
   END FE_OFN11522_n_140234

   PIN FE_OFN11557_n_137230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.186 0.0 51.214 0.163 ;
      END
   END FE_OFN11557_n_137230

   PIN FE_OFN11558_n_137230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.45 0.0 22.478 0.163 ;
      END
   END FE_OFN11558_n_137230

   PIN FE_OFN11607_n_39244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.45 0.0 70.478 0.163 ;
      END
   END FE_OFN11607_n_39244

   PIN FE_OFN11703_n_36821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.962 0.0 54.99 0.163 ;
      END
   END FE_OFN11703_n_36821

   PIN FE_OFN11879_n_143202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.29 0.0 74.318 0.163 ;
      END
   END FE_OFN11879_n_143202

   PIN FE_OFN11932_n_142850
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.114 0.0 96.142 0.163 ;
      END
   END FE_OFN11932_n_142850

   PIN FE_OFN12024_n_41611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.634 249.792 11.662 ;
      END
   END FE_OFN12024_n_41611

   PIN FE_OFN12028_n_143507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.458 0.0 73.486 0.163 ;
      END
   END FE_OFN12028_n_143507

   PIN FE_OFN12037_n_143629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.514 249.792 38.542 ;
      END
   END FE_OFN12037_n_143629

   PIN FE_OFN12040_n_143629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.386 0.0 246.414 0.163 ;
      END
   END FE_OFN12040_n_143629

   PIN FE_OFN12061_n_143423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.154 249.792 55.182 ;
      END
   END FE_OFN12061_n_143423

   PIN FE_OFN12085_n_143619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.33 0.0 97.358 0.163 ;
      END
   END FE_OFN12085_n_143619

   PIN FE_OFN12624_n_143670
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.586 249.792 49.614 ;
      END
   END FE_OFN12624_n_143670

   PIN FE_OFN12632_n_143496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.418 249.792 18.446 ;
      END
   END FE_OFN12632_n_143496

   PIN FE_OFN12753_n_142961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.162 0.0 50.19 0.163 ;
      END
   END FE_OFN12753_n_142961

   PIN FE_OFN12761_n_41012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.354 249.792 18.382 ;
      END
   END FE_OFN12761_n_41012

   PIN FE_OFN12764_n_41015
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.61 249.792 26.638 ;
      END
   END FE_OFN12764_n_41015

   PIN FE_OFN12968_n_112030
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.994 0.0 51.022 0.163 ;
      END
   END FE_OFN12968_n_112030

   PIN FE_OFN13044_n_40829
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.266 249.792 57.294 ;
      END
   END FE_OFN13044_n_40829

   PIN FE_OFN13226_n_143481
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.41 249.792 15.438 ;
      END
   END FE_OFN13226_n_143481

   PIN FE_OFN13233_n_143479
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.01 249.792 41.038 ;
      END
   END FE_OFN13233_n_143479

   PIN FE_OFN13239_n_41374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 47.602 249.792 47.63 ;
      END
   END FE_OFN13239_n_41374

   PIN FE_OFN13242_n_41374
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.81 249.792 45.838 ;
      END
   END FE_OFN13242_n_41374

   PIN FE_OFN13246_n_143370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 46.066 249.792 46.094 ;
      END
   END FE_OFN13246_n_143370

   PIN FE_OFN13253_n_143369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.946 249.792 40.974 ;
      END
   END FE_OFN13253_n_143369

   PIN FE_OFN13297_n_143032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.386 0.0 70.414 0.163 ;
      END
   END FE_OFN13297_n_143032

   PIN FE_OFN13347_n_142796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.442 0.0 43.47 0.163 ;
      END
   END FE_OFN13347_n_142796

   PIN FE_OFN13348_n_142796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.994 0.0 59.022 0.163 ;
      END
   END FE_OFN13348_n_142796

   PIN FE_OFN13393_n_41612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 23.346 249.792 23.374 ;
      END
   END FE_OFN13393_n_41612

   PIN FE_OFN13450_n_41900
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.45 249.792 62.478 ;
      END
   END FE_OFN13450_n_41900

   PIN FE_OFN13460_n_42034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 91.954 249.792 91.982 ;
      END
   END FE_OFN13460_n_42034

   PIN FE_OFN13515_n_112357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.866 0.0 34.894 0.163 ;
      END
   END FE_OFN13515_n_112357

   PIN FE_OFN13525_n_137232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.314 0.0 51.342 0.163 ;
      END
   END FE_OFN13525_n_137232

   PIN FE_OFN13528_n_137233
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.346 249.792 15.374 ;
      END
   END FE_OFN13528_n_137233

   PIN FE_OFN13529_n_137233
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.194 249.792 30.222 ;
      END
   END FE_OFN13529_n_137233

   PIN FE_OFN13672_n_143509
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.402 0.0 52.43 0.163 ;
      END
   END FE_OFN13672_n_143509

   PIN FE_OFN13686_n_143426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 19.058 249.792 19.086 ;
      END
   END FE_OFN13686_n_143426

   PIN FE_OFN13777_n_41686
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.09 0.0 55.118 0.163 ;
      END
   END FE_OFN13777_n_41686

   PIN FE_OFN13787_n_41960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 4.018 249.792 4.046 ;
      END
   END FE_OFN13787_n_41960

   PIN FE_OFN13789_n_41995
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 13.682 249.792 13.71 ;
      END
   END FE_OFN13789_n_41995

   PIN FE_OFN13796_n_41995
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.834 249.792 30.862 ;
      END
   END FE_OFN13796_n_41995

   PIN FE_OFN13864_n_41964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 40.626 249.792 40.654 ;
      END
   END FE_OFN13864_n_41964

   PIN FE_OFN14082_n_142962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.69 0.0 64.718 0.163 ;
      END
   END FE_OFN14082_n_142962

   PIN FE_OFN14361_n_143300
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.194 0.0 78.222 0.082 ;
      END
   END FE_OFN14361_n_143300

   PIN FE_OFN14401_n_142794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.162 0.0 90.19 0.163 ;
      END
   END FE_OFN14401_n_142794

   PIN FE_OFN14406_n_31761
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.802 0.0 58.83 0.163 ;
      END
   END FE_OFN14406_n_31761

   PIN FE_OFN14899_n_140203
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.882 249.792 40.91 ;
      END
   END FE_OFN14899_n_140203

   PIN FE_OFN15134_n_30145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 58.29 249.792 58.318 ;
      END
   END FE_OFN15134_n_30145

   PIN FE_OFN15168_n_31480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 111.602 249.792 111.63 ;
      END
   END FE_OFN15168_n_31480

   PIN FE_OFN15328_n_29953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 248.882 0.0 248.91 0.163 ;
      END
   END FE_OFN15328_n_29953

   PIN FE_OFN15342_n_30559
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.698 0.0 235.726 0.163 ;
      END
   END FE_OFN15342_n_30559

   PIN FE_OFN16113_n_42033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 69.106 249.792 69.134 ;
      END
   END FE_OFN16113_n_42033

   PIN FE_OFN17005_n_58282
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 212.594 117.597 212.622 117.76 ;
      END
   END FE_OFN17005_n_58282

   PIN FE_OFN17026_n_66756
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 231.858 117.597 231.886 117.76 ;
      END
   END FE_OFN17026_n_66756

   PIN FE_OFN17099_n_53555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.802 249.792 106.83 ;
      END
   END FE_OFN17099_n_53555

   PIN FE_OFN17825_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.978 249.792 85.006 ;
      END
   END FE_OFN17825_delay_mul_ln34_unr7_unr0_stage2_stallmux_z_12_

   PIN FE_OFN17835_n_84330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.458 249.792 49.486 ;
      END
   END FE_OFN17835_n_84330

   PIN FE_OFN17869_n_65432
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.906 249.792 57.934 ;
      END
   END FE_OFN17869_n_65432

   PIN FE_OFN17921_n_57488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.738 249.792 18.766 ;
      END
   END FE_OFN17921_n_57488

   PIN FE_OFN17931_n_41611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.218 249.792 55.246 ;
      END
   END FE_OFN17931_n_41611

   PIN FE_OFN18301_b_4_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.666 0.0 47.694 0.163 ;
      END
   END FE_OFN18301_b_4_4_4

   PIN FE_OFN18306_b_4_8_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 73.586 0.0 73.614 0.163 ;
      END
   END FE_OFN18306_b_4_8_5

   PIN FE_OFN18401_n_31516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.746 249.792 45.774 ;
      END
   END FE_OFN18401_n_31516

   PIN FE_OFN18434_n_27857
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.498 0.0 216.526 0.163 ;
      END
   END FE_OFN18434_n_27857

   PIN FE_OFN18783_n_31306
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 96.05 249.792 96.078 ;
      END
   END FE_OFN18783_n_31306

   PIN FE_OFN18962_n_41993
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.57 249.792 11.598 ;
      END
   END FE_OFN18962_n_41993

   PIN FE_OFN18995_n_41993
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 61.106 249.792 61.134 ;
      END
   END FE_OFN18995_n_41993

   PIN FE_OFN2320_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.906 117.597 241.934 117.76 ;
      END
   END FE_OFN2320_delay_mul_ln34_unr9_unr7_stage2_stallmux_z_14_

   PIN FE_OFN4455_n_10397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.914 0.0 12.942 0.163 ;
      END
   END FE_OFN4455_n_10397

   PIN FE_OFN4458_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.098 0.0 18.126 0.163 ;
      END
   END FE_OFN4458_delay_mul_ln34_unr4_unr2_stage2_stallmux_z_12_

   PIN FE_OFN4574_n_142961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.426 0.0 37.454 0.163 ;
      END
   END FE_OFN4574_n_142961

   PIN FE_OFN4623_n_142793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.346 0.0 47.374 0.082 ;
      END
   END FE_OFN4623_n_142793

   PIN FE_OFN4667_n_137232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.562 0.0 24.59 0.163 ;
      END
   END FE_OFN4667_n_137232

   PIN FE_OFN4683_n_143620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.026 0.0 79.054 0.163 ;
      END
   END FE_OFN4683_n_143620

   PIN FE_OFN4730_n_143033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.058 0.0 83.086 0.163 ;
      END
   END FE_OFN4730_n_143033

   PIN FE_OFN4781_n_143003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.962 0.0 38.99 0.163 ;
      END
   END FE_OFN4781_n_143003

   PIN FE_OFN4821_n_143199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.954 0.0 35.982 0.163 ;
      END
   END FE_OFN4821_n_143199

   PIN FE_OFN4837_n_140222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.378 0.0 51.406 0.163 ;
      END
   END FE_OFN4837_n_140222

   PIN FE_OFN4869_n_143507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.922 0.0 31.95 0.163 ;
      END
   END FE_OFN4869_n_143507

   PIN FE_OFN4891_n_140207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 56.562 0.0 56.59 0.163 ;
      END
   END FE_OFN4891_n_140207

   PIN FE_OFN6426_n_45151
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.322 249.792 62.35 ;
      END
   END FE_OFN6426_n_45151

   PIN FE_OFN6603_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 48.754 249.792 48.782 ;
      END
   END FE_OFN6603_n_140234

   PIN FE_OFN6604_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 38.386 249.792 38.414 ;
      END
   END FE_OFN6604_n_140234

   PIN FE_OFN6610_n_140234
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 25.97 249.792 25.998 ;
      END
   END FE_OFN6610_n_140234

   PIN FE_OFN6660_n_41611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.01 249.792 33.038 ;
      END
   END FE_OFN6660_n_41611

   PIN FE_OFN6723_n_41706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.586 249.792 57.614 ;
      END
   END FE_OFN6723_n_41706

   PIN FE_OFN6734_n_41994
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.202 249.792 57.23 ;
      END
   END FE_OFN6734_n_41994

   PIN FE_OFN6770_n_143423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.818 249.792 40.846 ;
      END
   END FE_OFN6770_n_143423

   PIN FE_OFN6842_n_41015
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.538 249.792 55.566 ;
      END
   END FE_OFN6842_n_41015

   PIN FE_OFN6876_n_41734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.71 65.266 249.792 65.294 ;
      END
   END FE_OFN6876_n_41734

   PIN FE_OFN6961_n_140210
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.41 249.792 55.438 ;
      END
   END FE_OFN6961_n_140210

   PIN FE_OFN7004_n_140202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 40.562 249.792 40.59 ;
      END
   END FE_OFN7004_n_140202

   PIN FE_OFN7022_n_66979
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.642 249.792 70.67 ;
      END
   END FE_OFN7022_n_66979

   PIN FE_OFN8169_n_26637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.954 117.597 227.982 117.76 ;
      END
   END FE_OFN8169_n_26637

   PIN FE_OFN8329_n_31307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 88.37 249.792 88.398 ;
      END
   END FE_OFN8329_n_31307

   PIN FE_OFN8463_n_25371
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 63.026 249.792 63.054 ;
      END
   END FE_OFN8463_n_25371

   PIN FE_OFN8477_n_30279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.538 0.0 239.566 0.163 ;
      END
   END FE_OFN8477_n_30279

   PIN FE_OFN8491_n_29557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 243.378 0.0 243.406 0.163 ;
      END
   END FE_OFN8491_n_29557

   PIN FE_OFN8577_n_29968
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.874 0.0 245.902 0.163 ;
      END
   END FE_OFN8577_n_29968

   PIN FE_OFN8703_n_31118
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.93 249.792 18.958 ;
      END
   END FE_OFN8703_n_31118

   PIN FE_OFN8799_n_25382
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.634 0.0 235.662 0.163 ;
      END
   END FE_OFN8799_n_25382

   PIN FE_OFN9238_delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.426 0.0 197.454 0.163 ;
      END
   END FE_OFN9238_delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_

   PIN FE_OFN9464_b_7_8_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 31.346 249.792 31.374 ;
      END
   END FE_OFN9464_b_7_8_11

   PIN FE_OFN9467_b_7_8_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.25 249.792 11.278 ;
      END
   END FE_OFN9467_b_7_8_10

   PIN FE_OFN9480_b_7_8_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.514 249.792 22.542 ;
      END
   END FE_OFN9480_b_7_8_5

   PIN FE_OFN9486_b_7_8_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 25.842 249.792 25.87 ;
      END
   END FE_OFN9486_b_7_8_3

   PIN FE_OFN9489_b_7_8_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.45 249.792 22.478 ;
      END
   END FE_OFN9489_b_7_8_2

   PIN FE_OFN9557_b_7_6_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.474 249.792 55.502 ;
      END
   END FE_OFN9557_b_7_6_6

   PIN FE_OFN9563_b_7_6_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 85.554 249.792 85.582 ;
      END
   END FE_OFN9563_b_7_6_5

   PIN FE_OFN9566_b_7_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.778 249.792 41.806 ;
      END
   END FE_OFN9566_b_7_6_4

   PIN FE_OFN9568_b_7_6_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 41.202 249.792 41.23 ;
      END
   END FE_OFN9568_b_7_6_3

   PIN FE_OFN9573_b_7_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 61.234 249.792 61.262 ;
      END
   END FE_OFN9573_b_7_6_2

   PIN FE_OFN9575_b_7_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.002 249.792 38.03 ;
      END
   END FE_OFN9575_b_7_6_2

   PIN FE_OFN9576_b_7_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.338 117.597 220.366 117.76 ;
      END
   END FE_OFN9576_b_7_6_1

   PIN FE_OFN9580_b_7_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.71 34.034 249.792 34.062 ;
      END
   END FE_OFN9580_b_7_6_0

   PIN FE_OFN9732_b_7_0_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 64.882 249.792 64.91 ;
      END
   END FE_OFN9732_b_7_0_10

   PIN FE_OFN9735_b_7_0_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 55.346 249.792 55.374 ;
      END
   END FE_OFN9735_b_7_0_9

   PIN FE_OFN9752_b_7_0_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.002 249.792 70.03 ;
      END
   END FE_OFN9752_b_7_0_5

   PIN FE_OFN9757_b_7_0_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.386 249.792 62.414 ;
      END
   END FE_OFN9757_b_7_0_4

   PIN FE_OFN9765_b_7_0_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.71 62.77 249.792 62.798 ;
      END
   END FE_OFN9765_b_7_0_2

   PIN FE_OFN9769_b_7_0_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 49.778 249.792 49.806 ;
      END
   END FE_OFN9769_b_7_0_1

   PIN FE_OFN9772_b_7_0_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 72.946 249.792 72.974 ;
      END
   END FE_OFN9772_b_7_0_0

   PIN FE_OFN9858_b_4_8_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.682 0.0 61.71 0.163 ;
      END
   END FE_OFN9858_b_4_8_13

   PIN FE_OFN9860_b_4_8_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.834 0.0 62.862 0.163 ;
      END
   END FE_OFN9860_b_4_8_12

   PIN FE_OFN9862_b_4_8_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.77 0.0 62.798 0.163 ;
      END
   END FE_OFN9862_b_4_8_11

   PIN FE_OFN9883_b_4_8_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 70.514 0.0 70.542 0.082 ;
      END
   END FE_OFN9883_b_4_8_2

   PIN FE_OFN9961_b_4_6_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.09 0.0 79.118 0.082 ;
      END
   END FE_OFN9961_b_4_6_3

   PIN FE_OFN9964_b_4_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.762 0.0 75.79 0.082 ;
      END
   END FE_OFN9964_b_4_6_2

   PIN b_4_8_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.266 117.597 105.294 117.76 ;
      END
   END b_4_8_3

   PIN b_7_0_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 72.882 249.792 72.91 ;
      END
   END b_7_0_7

   PIN b_7_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 55.282 249.792 55.31 ;
      END
   END b_7_6_0

   PIN b_7_6_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.978 117.597 205.006 117.76 ;
      END
   END b_7_6_10

   PIN b_7_6_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 206.45 117.597 206.478 117.76 ;
      END
   END b_7_6_11

   PIN b_7_6_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 220.402 117.597 220.43 117.76 ;
      END
   END b_7_6_14

   PIN b_7_6_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 216.818 117.597 216.846 117.76 ;
      END
   END b_7_6_15

   PIN b_7_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 229.49 117.597 229.518 117.76 ;
      END
   END b_7_6_4

   PIN b_7_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 62.962 249.792 62.99 ;
      END
   END b_7_6_7

   PIN b_7_6_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 220.338 117.597 220.366 117.76 ;
      END
   END b_7_6_9

   PIN b_7_8_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 171.762 117.597 171.79 117.76 ;
      END
   END b_7_8_7

   PIN b_7_8_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 197.298 117.597 197.326 117.76 ;
      END
   END b_7_8_8

   PIN delay_mul_ln34_unr7_unr8_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 174.642 0.0 174.67 0.163 ;
      END
   END delay_mul_ln34_unr7_unr8_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr8_unr1_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.57 249.792 99.598 ;
      END
   END delay_mul_ln34_unr8_unr1_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr8_unr7_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.946 249.792 32.974 ;
      END
   END delay_mul_ln34_unr8_unr7_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr8_unr7_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 18.226 249.792 18.254 ;
      END
   END delay_mul_ln34_unr8_unr7_stage2_stallmux_z_3_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.658 117.597 212.686 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.466 117.597 220.494 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr9_unr7_stage2_stallmux_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.498 117.597 216.526 117.76 ;
      END
   END delay_mul_ln34_unr9_unr7_stage2_stallmux_z_3_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.802 117.678 66.83 117.76 ;
      END
   END ispd_clk

   PIN mul_4647_72_n_181
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.298 0.0 5.326 0.163 ;
      END
   END mul_4647_72_n_181

   PIN mul_4647_72_n_182
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.69 0.0 16.718 0.163 ;
      END
   END mul_4647_72_n_182

   PIN mul_4647_72_n_53
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.426 0.0 5.454 0.163 ;
      END
   END mul_4647_72_n_53

   PIN mul_4647_72_n_69
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.154 0.0 7.182 0.163 ;
      END
   END mul_4647_72_n_69

   PIN mul_4647_72_n_779
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.562 0.163 40.59 ;
      END
   END mul_4647_72_n_779

   PIN mul_4649_72_n_825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.562 0.0 120.59 0.163 ;
      END
   END mul_4649_72_n_825

   PIN mul_4649_72_n_88
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.69 0.0 112.718 0.163 ;
      END
   END mul_4649_72_n_88

   PIN mul_4651_72_n_285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.386 0.0 94.414 0.163 ;
      END
   END mul_4651_72_n_285

   PIN mul_4664_72_n_241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.738 0.0 74.766 0.163 ;
      END
   END mul_4664_72_n_241

   PIN mul_4664_72_n_242
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.25 0.0 75.278 0.163 ;
      END
   END mul_4664_72_n_242

   PIN mul_4664_72_n_317
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.818 0.0 56.846 0.163 ;
      END
   END mul_4664_72_n_317

   PIN mul_4664_72_n_318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.754 0.0 56.782 0.163 ;
      END
   END mul_4664_72_n_318

   PIN mul_4664_72_n_319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.386 0.0 54.414 0.163 ;
      END
   END mul_4664_72_n_319

   PIN mul_4664_72_n_813
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.882 0.0 32.91 0.163 ;
      END
   END mul_4664_72_n_813

   PIN mul_4664_72_n_825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.386 0.0 62.414 0.163 ;
      END
   END mul_4664_72_n_825

   PIN mul_4664_72_n_84
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.706 0.0 62.734 0.163 ;
      END
   END mul_4664_72_n_84

   PIN mul_4664_72_n_848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.562 0.0 32.59 0.163 ;
      END
   END mul_4664_72_n_848

   PIN mul_4664_72_n_85
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.474 0.0 71.502 0.163 ;
      END
   END mul_4664_72_n_85

   PIN mul_4664_72_n_88
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.714 0.0 41.742 0.163 ;
      END
   END mul_4664_72_n_88

   PIN mul_4698_72_n_100
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.602 249.792 7.63 ;
      END
   END mul_4698_72_n_100

   PIN mul_4698_72_n_99
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.89 249.792 3.918 ;
      END
   END mul_4698_72_n_99

   PIN mul_4700_72_n_178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 8.114 249.792 8.142 ;
      END
   END mul_4700_72_n_178

   PIN mul_4700_72_n_179
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.826 249.792 3.854 ;
      END
   END mul_4700_72_n_179

   PIN n_101492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.762 249.792 3.79 ;
      END
   END n_101492

   PIN n_102695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 193.138 117.597 193.166 117.76 ;
      END
   END n_102695

   PIN n_103071
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.626 117.597 216.654 117.76 ;
      END
   END n_103071

   PIN n_103939
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 225.522 117.597 225.55 117.76 ;
      END
   END n_103939

   PIN n_103940
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 232.562 117.597 232.59 117.76 ;
      END
   END n_103940

   PIN n_106720
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 114.226 249.792 114.254 ;
      END
   END n_106720

   PIN n_107989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.378 0.0 43.406 0.163 ;
      END
   END n_107989

   PIN n_108267
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.69 117.597 208.718 117.76 ;
      END
   END n_108267

   PIN n_108268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.89 117.597 203.918 117.76 ;
      END
   END n_108268

   PIN n_108688
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 189.554 117.597 189.582 117.76 ;
      END
   END n_108688

   PIN n_110443
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.434 249.792 80.462 ;
      END
   END n_110443

   PIN n_110533
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.074 117.597 201.102 117.76 ;
      END
   END n_110533

   PIN n_112122
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 84.722 0.163 84.75 ;
      END
   END n_112122

   PIN n_112183
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.09 0.0 63.118 0.082 ;
      END
   END n_112183

   PIN n_112413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.49 0.0 93.518 0.163 ;
      END
   END n_112413

   PIN n_112659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 75.186 0.0 75.214 0.163 ;
      END
   END n_112659

   PIN n_114178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.794 0.0 47.822 0.163 ;
      END
   END n_114178

   PIN n_114182
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.658 0.0 12.686 0.163 ;
      END
   END n_114182

   PIN n_114494
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.146 0.0 28.174 0.163 ;
      END
   END n_114494

   PIN n_114496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.082 0.0 28.11 0.163 ;
      END
   END n_114496

   PIN n_114524
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.722 0.0 12.75 0.163 ;
      END
   END n_114524

   PIN n_114615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.61 0.0 42.638 0.163 ;
      END
   END n_114615

   PIN n_114617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.114 0.0 24.142 0.163 ;
      END
   END n_114617

   PIN n_114672
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.754 117.597 48.782 117.76 ;
      END
   END n_114672

   PIN n_114673
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.21 0.0 28.238 0.163 ;
      END
   END n_114673

   PIN n_114676
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.05 0.0 24.078 0.163 ;
      END
   END n_114676

   PIN n_114855
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.954 0.0 43.982 0.163 ;
      END
   END n_114855

   PIN n_114920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.93 0.0 58.958 0.163 ;
      END
   END n_114920

   PIN n_114921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 58.738 0.0 58.766 0.163 ;
      END
   END n_114921

   PIN n_115152
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.466 0.0 52.494 0.163 ;
      END
   END n_115152

   PIN n_115153
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.274 0.0 52.302 0.163 ;
      END
   END n_115153

   PIN n_115190
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.658 0.0 44.686 0.163 ;
      END
   END n_115190

   PIN n_115308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.05 0.0 32.078 0.163 ;
      END
   END n_115308

   PIN n_115309
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.21 0.0 28.238 0.163 ;
      END
   END n_115309

   PIN n_115311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.538 0.0 47.566 0.163 ;
      END
   END n_115311

   PIN n_115543
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.946 0.0 8.974 0.163 ;
      END
   END n_115543

   PIN n_115582
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.698 0.0 35.726 0.163 ;
      END
   END n_115582

   PIN n_115593
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.85 0.0 20.878 0.163 ;
      END
   END n_115593

   PIN n_115606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.698 0.0 43.726 0.163 ;
      END
   END n_115606

   PIN n_115661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.57 0.0 51.598 0.163 ;
      END
   END n_115661

   PIN n_115793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.602 0.0 47.63 0.163 ;
      END
   END n_115793

   PIN n_115794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.474 0.0 47.502 0.163 ;
      END
   END n_115794

   PIN n_115810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.562 0.0 16.59 0.163 ;
      END
   END n_115810

   PIN n_116281
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.73 0.0 39.758 0.163 ;
      END
   END n_116281

   PIN n_116796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.93 0.0 34.958 0.163 ;
      END
   END n_116796

   PIN n_117132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.786 0.0 76.814 0.163 ;
      END
   END n_117132

   PIN n_117734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.242 0.0 24.27 0.163 ;
      END
   END n_117734

   PIN n_117835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.826 0.0 35.854 0.163 ;
      END
   END n_117835

   PIN n_118212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.41 0.0 47.438 0.163 ;
      END
   END n_118212

   PIN n_118398
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.178 0.0 16.206 0.163 ;
      END
   END n_118398

   PIN n_119074
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.162 0.163 114.19 ;
      END
   END n_119074

   PIN n_120882
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.634 117.597 43.662 117.76 ;
      END
   END n_120882

   PIN n_121314
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.274 0.0 28.302 0.163 ;
      END
   END n_121314

   PIN n_121751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.114 0.0 32.142 0.163 ;
      END
   END n_121751

   PIN n_121989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.37 0.0 24.398 0.163 ;
      END
   END n_121989

   PIN n_122315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.178 0.0 24.206 0.163 ;
      END
   END n_122315

   PIN n_122349
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.634 0.0 35.662 0.163 ;
      END
   END n_122349

   PIN n_123446
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.218 0.0 47.246 0.163 ;
      END
   END n_123446

   PIN n_124498
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.602 0.163 7.63 ;
      END
   END n_124498

   PIN n_124539
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.746 117.597 37.774 117.76 ;
      END
   END n_124539

   PIN n_124540
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.01 117.597 41.038 117.76 ;
      END
   END n_124540

   PIN n_124638
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.626 0.0 16.654 0.163 ;
      END
   END n_124638

   PIN n_124639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 24.562 0.0 24.59 0.163 ;
      END
   END n_124639

   PIN n_125192
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.626 117.597 8.654 117.76 ;
      END
   END n_125192

   PIN n_125461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.69 0.0 24.718 0.163 ;
      END
   END n_125461

   PIN n_125695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.938 0.0 21.966 0.163 ;
      END
   END n_125695

   PIN n_125716
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.618 0.0 13.646 0.163 ;
      END
   END n_125716

   PIN n_127036
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 12.85 0.0 12.878 0.163 ;
      END
   END n_127036

   PIN n_127040
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.002 0.0 30.03 0.163 ;
      END
   END n_127040

   PIN n_127190
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.05 117.597 48.078 117.76 ;
      END
   END n_127190

   PIN n_127195
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.746 0.0 13.774 0.163 ;
      END
   END n_127195

   PIN n_127589
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.466 0.163 4.494 ;
      END
   END n_127589

   PIN n_127666
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.818 117.597 24.846 117.76 ;
      END
   END n_127666

   PIN n_128129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.338 0.0 28.366 0.163 ;
      END
   END n_128129

   PIN n_128287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.506 0.0 3.534 0.163 ;
      END
   END n_128287

   PIN n_128296
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.202 0.0 9.23 0.163 ;
      END
   END n_128296

   PIN n_128768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.074 117.597 57.102 117.76 ;
      END
   END n_128768

   PIN n_129724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.33 0.0 9.358 0.163 ;
      END
   END n_129724

   PIN n_130012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.402 0.0 20.43 0.163 ;
      END
   END n_130012

   PIN n_130016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.498 0.0 16.526 0.163 ;
      END
   END n_130016

   PIN n_131230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.338 0.0 20.366 0.163 ;
      END
   END n_131230

   PIN n_132777
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.274 117.597 28.302 117.76 ;
      END
   END n_132777

   PIN n_133344
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.882 0.0 16.91 0.163 ;
      END
   END n_133344

   PIN n_133767
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.762 0.0 35.79 0.163 ;
      END
   END n_133767

   PIN n_137225
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.474 0.0 47.502 0.163 ;
      END
   END n_137225

   PIN n_137233
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.506 249.792 11.534 ;
      END
   END n_137233

   PIN n_137728
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.698 249.792 3.726 ;
      END
   END n_137728

   PIN n_137826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 34.162 249.792 34.19 ;
      END
   END n_137826

   PIN n_137827
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.906 0.0 65.934 0.163 ;
      END
   END n_137827

   PIN n_137828
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 89.778 0.0 89.806 0.163 ;
      END
   END n_137828

   PIN n_137851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.506 0.0 43.534 0.163 ;
      END
   END n_137851

   PIN n_140213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.386 249.792 70.414 ;
      END
   END n_140213

   PIN n_142851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.442 0.0 67.47 0.082 ;
      END
   END n_142851

   PIN n_142964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.546 0.0 66.574 0.163 ;
      END
   END n_142964

   PIN n_143483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.71 26.93 249.792 26.958 ;
      END
   END n_143483

   PIN n_143496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 27.186 249.792 27.214 ;
      END
   END n_143496

   PIN n_143630
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.682 249.792 45.71 ;
      END
   END n_143630

   PIN n_143743
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.554 0.0 13.582 0.163 ;
      END
   END n_143743

   PIN n_143933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.386 0.0 110.414 0.163 ;
      END
   END n_143933

   PIN n_144109
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.538 0.0 87.566 0.163 ;
      END
   END n_144109

   PIN n_144135
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.05 117.597 224.078 117.76 ;
      END
   END n_144135

   PIN n_144158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.474 249.792 47.502 ;
      END
   END n_144158

   PIN n_24056
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.442 249.792 3.47 ;
      END
   END n_24056

   PIN n_25134
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 171.25 0.0 171.278 0.163 ;
      END
   END n_25134

   PIN n_25376
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.618 249.792 45.646 ;
      END
   END n_25376

   PIN n_26011
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.386 0.0 166.414 0.163 ;
      END
   END n_26011

   PIN n_26383
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.25 117.597 147.278 117.76 ;
      END
   END n_26383

   PIN n_26633
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.738 249.792 106.766 ;
      END
   END n_26633

   PIN n_27338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 158.706 117.597 158.734 117.76 ;
      END
   END n_27338

   PIN n_27740
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.898 249.792 38.926 ;
      END
   END n_27740

   PIN n_27741
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.834 249.792 38.862 ;
      END
   END n_27741

   PIN n_28380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 4.53 249.792 4.558 ;
      END
   END n_28380

   PIN n_28496
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.946 117.597 208.974 117.76 ;
      END
   END n_28496

   PIN n_28631
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 124.338 0.0 124.366 0.163 ;
      END
   END n_28631

   PIN n_28640
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 4.466 249.792 4.494 ;
      END
   END n_28640

   PIN n_28780
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 208.882 117.597 208.91 117.76 ;
      END
   END n_28780

   PIN n_29125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 213.106 0.0 213.134 0.163 ;
      END
   END n_29125

   PIN n_31876
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.85 0.0 92.878 0.163 ;
      END
   END n_31876

   PIN n_33226
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.154 0.0 47.182 0.163 ;
      END
   END n_33226

   PIN n_33292
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.746 0.0 85.774 0.163 ;
      END
   END n_33292

   PIN n_33293
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.402 0.0 84.43 0.163 ;
      END
   END n_33293

   PIN n_33375
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.962 0.0 62.99 0.163 ;
      END
   END n_33375

   PIN n_33782
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.842 0.0 81.87 0.163 ;
      END
   END n_33782

   PIN n_34260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.562 249.792 40.59 ;
      END
   END n_34260

   PIN n_34345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.674 0.0 66.702 0.163 ;
      END
   END n_34345

   PIN n_35072
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.554 0.0 69.582 0.163 ;
      END
   END n_35072

   PIN n_35096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.786 0.0 116.814 0.163 ;
      END
   END n_35096

   PIN n_36000
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.49 0.0 69.518 0.163 ;
      END
   END n_36000

   PIN n_36612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.218 0.0 71.246 0.163 ;
      END
   END n_36612

   PIN n_37235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.45 0.0 54.478 0.163 ;
      END
   END n_37235

   PIN n_37476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.442 0.0 67.47 0.163 ;
      END
   END n_37476

   PIN n_40827
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 27.122 249.792 27.15 ;
      END
   END n_40827

   PIN n_40897
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.634 249.792 3.662 ;
      END
   END n_40897

   PIN n_40960
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 8.946 249.792 8.974 ;
      END
   END n_40960

   PIN n_41417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 23.282 249.792 23.31 ;
      END
   END n_41417

   PIN n_41500
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.57 249.792 3.598 ;
      END
   END n_41500

   PIN n_41612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.282 249.792 15.31 ;
      END
   END n_41612

   PIN n_41734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.77 249.792 30.798 ;
      END
   END n_41734

   PIN n_41834
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.922 249.792 7.95 ;
      END
   END n_41834

   PIN n_41962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 11.186 249.792 11.214 ;
      END
   END n_41962

   PIN n_42268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 78.002 249.792 78.03 ;
      END
   END n_42268

   PIN n_42269
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.938 249.792 77.966 ;
      END
   END n_42269

   PIN n_42354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.474 249.792 103.502 ;
      END
   END n_42354

   PIN n_42362
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 107.25 249.792 107.278 ;
      END
   END n_42362

   PIN n_42412
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.874 249.792 77.902 ;
      END
   END n_42412

   PIN n_42413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.81 249.792 77.838 ;
      END
   END n_42413

   PIN n_42443
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.546 249.792 106.574 ;
      END
   END n_42443

   PIN n_42504
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 88.178 249.792 88.206 ;
      END
   END n_42504

   PIN n_42506
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 95.922 249.792 95.95 ;
      END
   END n_42506

   PIN n_42608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.482 249.792 106.51 ;
      END
   END n_42608

   PIN n_42807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 111.538 249.792 111.566 ;
      END
   END n_42807

   PIN n_42921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 243.378 117.597 243.406 117.76 ;
      END
   END n_42921

   PIN n_43096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.77 249.792 70.798 ;
      END
   END n_43096

   PIN n_43134
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.41 249.792 103.438 ;
      END
   END n_43134

   PIN n_43240
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.282 249.792 103.31 ;
      END
   END n_43240

   PIN n_43320
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.522 249.792 57.55 ;
      END
   END n_43320

   PIN n_43384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 114.354 249.792 114.382 ;
      END
   END n_43384

   PIN n_43416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 91.89 249.792 91.918 ;
      END
   END n_43416

   PIN n_43545
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.706 249.792 70.734 ;
      END
   END n_43545

   PIN n_43643
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 85.106 249.792 85.134 ;
      END
   END n_43643

   PIN n_43707
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 99.442 249.792 99.47 ;
      END
   END n_43707

   PIN n_44058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.346 249.792 103.374 ;
      END
   END n_44058

   PIN n_44137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.73 117.597 231.758 117.76 ;
      END
   END n_44137

   PIN n_44356
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.13 249.792 30.158 ;
      END
   END n_44356

   PIN n_44415
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.322 249.792 70.35 ;
      END
   END n_44415

   PIN n_44594
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 107.314 249.792 107.342 ;
      END
   END n_44594

   PIN n_44658
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 107.186 249.792 107.214 ;
      END
   END n_44658

   PIN n_45114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 111.346 249.792 111.374 ;
      END
   END n_45114

   PIN n_45130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.258 249.792 70.286 ;
      END
   END n_45130

   PIN n_45297
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.194 249.792 70.222 ;
      END
   END n_45297

   PIN n_45432
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.546 249.792 26.574 ;
      END
   END n_45432

   PIN n_45433
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 27.058 249.792 27.086 ;
      END
   END n_45433

   PIN n_45435
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 73.202 249.792 73.23 ;
      END
   END n_45435

   PIN n_45598
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 91.762 249.792 91.79 ;
      END
   END n_45598

   PIN n_45795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.914 249.792 84.942 ;
      END
   END n_45795

   PIN n_45796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.85 249.792 84.878 ;
      END
   END n_45796

   PIN n_46004
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 33.522 249.792 33.55 ;
      END
   END n_46004

   PIN n_46071
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 23.218 249.792 23.246 ;
      END
   END n_46071

   PIN n_46080
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 46.066 249.792 46.094 ;
      END
   END n_46080

   PIN n_46178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.514 0.0 86.542 0.163 ;
      END
   END n_46178

   PIN n_46181
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.866 249.792 26.894 ;
      END
   END n_46181

   PIN n_46217
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.13 249.792 70.158 ;
      END
   END n_46217

   PIN n_46227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.602 249.792 47.63 ;
      END
   END n_46227

   PIN n_46333
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.37 249.792 48.398 ;
      END
   END n_46333

   PIN n_46334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 248.946 0.0 248.974 0.163 ;
      END
   END n_46334

   PIN n_46340
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.482 249.792 26.51 ;
      END
   END n_46340

   PIN n_46341
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.418 249.792 26.446 ;
      END
   END n_46341

   PIN n_46365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.858 249.792 7.886 ;
      END
   END n_46365

   PIN n_46513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 23.154 249.792 23.182 ;
      END
   END n_46513

   PIN n_46588
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 40.754 249.792 40.782 ;
      END
   END n_46588

   PIN n_46658
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.186 249.792 11.214 ;
      END
   END n_46658

   PIN n_46660
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.602 249.792 15.63 ;
      END
   END n_46660

   PIN n_46774
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 3.506 249.792 3.534 ;
      END
   END n_46774

   PIN n_46851
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 31.218 249.792 31.246 ;
      END
   END n_46851

   PIN n_46932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 37.938 249.792 37.966 ;
      END
   END n_46932

   PIN n_46954
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 19.058 249.792 19.086 ;
      END
   END n_46954

   PIN n_47028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.354 249.792 26.382 ;
      END
   END n_47028

   PIN n_47607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.442 0.0 51.47 0.163 ;
      END
   END n_47607

   PIN n_47644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.794 249.792 7.822 ;
      END
   END n_47644

   PIN n_47750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.89 0.0 83.918 0.163 ;
      END
   END n_47750

   PIN n_47929
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.594 0.0 60.622 0.163 ;
      END
   END n_47929

   PIN n_48546
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 38.962 249.792 38.99 ;
      END
   END n_48546

   PIN n_48611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.914 0.0 44.942 0.163 ;
      END
   END n_48611

   PIN n_48880
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 63.09 249.792 63.118 ;
      END
   END n_48880

   PIN n_48997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 19.186 249.792 19.214 ;
      END
   END n_48997

   PIN n_49055
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 23.026 249.792 23.054 ;
      END
   END n_49055

   PIN n_49568
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.138 0.0 9.166 0.163 ;
      END
   END n_49568

   PIN n_49769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.73 249.792 7.758 ;
      END
   END n_49769

   PIN n_49987
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.066 249.792 70.094 ;
      END
   END n_49987

   PIN n_50107
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 7.666 249.792 7.694 ;
      END
   END n_50107

   PIN n_50238
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 111.282 249.792 111.31 ;
      END
   END n_50238

   PIN n_50246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 81.01 249.792 81.038 ;
      END
   END n_50246

   PIN n_50397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.642 249.792 62.67 ;
      END
   END n_50397

   PIN n_50495
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 111.474 249.792 111.502 ;
      END
   END n_50495

   PIN n_50522
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.618 117.597 229.646 117.76 ;
      END
   END n_50522

   PIN n_50818
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 91.826 249.792 91.854 ;
      END
   END n_50818

   PIN n_50937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.73 0.0 191.758 0.163 ;
      END
   END n_50937

   PIN n_51078
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.394 249.792 65.422 ;
      END
   END n_51078

   PIN n_51110
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.29 249.792 26.318 ;
      END
   END n_51110

   PIN n_51111
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.226 249.792 26.254 ;
      END
   END n_51111

   PIN n_51211
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.706 249.792 30.734 ;
      END
   END n_51211

   PIN n_51212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 32.946 249.792 32.974 ;
      END
   END n_51212

   PIN n_51988
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.578 249.792 70.606 ;
      END
   END n_51988

   PIN n_52066
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.666 0.0 191.694 0.163 ;
      END
   END n_52066

   PIN n_52279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.674 249.792 106.702 ;
      END
   END n_52279

   PIN n_52455
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.498 249.792 80.526 ;
      END
   END n_52455

   PIN n_52456
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.37 249.792 80.398 ;
      END
   END n_52456

   PIN n_52502
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 32.882 249.792 32.91 ;
      END
   END n_52502

   PIN n_52697
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 111.41 249.792 111.438 ;
      END
   END n_52697

   PIN n_52749
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.538 249.792 103.566 ;
      END
   END n_52749

   PIN n_52750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.986 249.792 104.014 ;
      END
   END n_52750

   PIN n_52873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 95.73 249.792 95.758 ;
      END
   END n_52873

   PIN n_52994
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.138 249.792 57.166 ;
      END
   END n_52994

   PIN n_53090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 11.25 249.792 11.278 ;
      END
   END n_53090

   PIN n_53725
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.794 249.792 103.822 ;
      END
   END n_53725

   PIN n_53750
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.538 117.597 239.566 117.76 ;
      END
   END n_53750

   PIN n_53835
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.858 0.0 39.886 0.163 ;
      END
   END n_53835

   PIN n_54049
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 23.09 249.792 23.118 ;
      END
   END n_54049

   PIN n_54060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.666 249.792 15.694 ;
      END
   END n_54060

   PIN n_54354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 14.898 249.792 14.926 ;
      END
   END n_54354

   PIN n_54357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 11.122 249.792 11.15 ;
      END
   END n_54357

   PIN n_54358
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.442 249.792 11.47 ;
      END
   END n_54358

   PIN n_54853
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 53.746 249.792 53.774 ;
      END
   END n_54853

   PIN n_54873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 111.986 249.792 112.014 ;
      END
   END n_54873

   PIN n_54905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.474 117.597 239.502 117.76 ;
      END
   END n_54905

   PIN n_54906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.794 117.597 239.822 117.76 ;
      END
   END n_54906

   PIN n_54932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.666 117.597 231.694 117.76 ;
      END
   END n_54932

   PIN n_54940
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 107.506 249.792 107.534 ;
      END
   END n_54940

   PIN n_54943
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.306 117.597 216.334 117.76 ;
      END
   END n_54943

   PIN n_54953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.506 249.792 99.534 ;
      END
   END n_54953

   PIN n_55031
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 63.026 249.792 63.054 ;
      END
   END n_55031

   PIN n_55096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 19.122 249.792 19.15 ;
      END
   END n_55096

   PIN n_55097
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 26.162 249.792 26.19 ;
      END
   END n_55097

   PIN n_5512
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.722 0.0 20.75 0.163 ;
      END
   END n_5512

   PIN n_55141
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.57 117.597 235.598 117.76 ;
      END
   END n_55141

   PIN n_55158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.578 249.792 62.606 ;
      END
   END n_55158

   PIN n_55332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 95.922 249.792 95.95 ;
      END
   END n_55332

   PIN n_55444
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 23.026 249.792 23.054 ;
      END
   END n_55444

   PIN n_55445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 22.962 249.792 22.99 ;
      END
   END n_55445

   PIN n_55540
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.122 0.0 147.15 0.163 ;
      END
   END n_55540

   PIN n_55560
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 83.954 249.792 83.982 ;
      END
   END n_55560

   PIN n_55599
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 30.642 249.792 30.67 ;
      END
   END n_55599

   PIN n_55648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.058 0.0 147.086 0.163 ;
      END
   END n_55648

   PIN n_55722
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.21 0.0 140.238 0.163 ;
      END
   END n_55722

   PIN n_55790
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.89 249.792 11.918 ;
      END
   END n_55790

   PIN n_5584
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.674 0.0 10.702 0.163 ;
      END
   END n_5584

   PIN n_55908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 19.314 249.792 19.342 ;
      END
   END n_55908

   PIN n_56447
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 243.378 117.597 243.406 117.76 ;
      END
   END n_56447

   PIN n_56448
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 114.29 249.792 114.318 ;
      END
   END n_56448

   PIN n_56512
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.33 249.792 65.358 ;
      END
   END n_56512

   PIN n_56516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.266 249.792 65.294 ;
      END
   END n_56516

   PIN n_56956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 187.826 0.0 187.854 0.163 ;
      END
   END n_56956

   PIN n_57348
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 31.154 249.792 31.182 ;
      END
   END n_57348

   PIN n_57368
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 8.37 249.792 8.398 ;
      END
   END n_57368

   PIN n_57417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 31.09 249.792 31.118 ;
      END
   END n_57417

   PIN n_57444
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.858 0.0 231.886 0.163 ;
      END
   END n_57444

   PIN n_57615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.73 117.597 239.758 117.76 ;
      END
   END n_57615

   PIN n_57620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.218 0.0 55.246 0.163 ;
      END
   END n_57620

   PIN n_57624
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 77.106 249.792 77.134 ;
      END
   END n_57624

   PIN n_57629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 48.306 249.792 48.334 ;
      END
   END n_57629

   PIN n_57726
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 57.97 249.792 57.998 ;
      END
   END n_57726

   PIN n_57746
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.754 249.792 40.782 ;
      END
   END n_57746

   PIN n_57903
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.202 117.597 113.23 117.76 ;
      END
   END n_57903

   PIN n_57935
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.458 249.792 65.486 ;
      END
   END n_57935

   PIN n_57983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 163.89 117.597 163.918 117.76 ;
      END
   END n_57983

   PIN n_58082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 106.61 249.792 106.638 ;
      END
   END n_58082

   PIN n_58177
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 111.666 249.792 111.694 ;
      END
   END n_58177

   PIN n_58261
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.242 117.597 216.27 117.76 ;
      END
   END n_58261

   PIN n_58290
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 217.074 117.597 217.102 117.76 ;
      END
   END n_58290

   PIN n_58294
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 217.01 117.597 217.038 117.76 ;
      END
   END n_58294

   PIN n_58385
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 22.962 249.792 22.99 ;
      END
   END n_58385

   PIN n_58399
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.29 249.792 18.318 ;
      END
   END n_58399

   PIN n_58400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.226 249.792 18.254 ;
      END
   END n_58400

   PIN n_58672
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 65.586 249.792 65.614 ;
      END
   END n_58672

   PIN n_58674
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 15.218 249.792 15.246 ;
      END
   END n_58674

   PIN n_59053
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.538 249.792 47.566 ;
      END
   END n_59053

   PIN n_59056
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 73.138 249.792 73.166 ;
      END
   END n_59056

   PIN n_59131
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 18.162 249.792 18.19 ;
      END
   END n_59131

   PIN n_59166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.506 117.597 235.534 117.76 ;
      END
   END n_59166

   PIN n_59286
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.89 117.597 227.918 117.76 ;
      END
   END n_59286

   PIN n_59394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.402 117.597 220.43 117.76 ;
      END
   END n_59394

   PIN n_59605
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.25 0.0 147.278 0.163 ;
      END
   END n_59605

   PIN n_60089
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.666 117.597 135.694 117.76 ;
      END
   END n_60089

   PIN n_60346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 61.042 249.792 61.07 ;
      END
   END n_60346

   PIN n_60369
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.594 0.0 212.622 0.163 ;
      END
   END n_60369

   PIN n_60370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.658 0.0 212.686 0.163 ;
      END
   END n_60370

   PIN n_60378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 72.754 249.792 72.782 ;
      END
   END n_60378

   PIN n_60427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.826 249.792 11.854 ;
      END
   END n_60427

   PIN n_60554
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 40.69 249.792 40.718 ;
      END
   END n_60554

   PIN n_60615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 45.554 249.792 45.582 ;
      END
   END n_60615

   PIN n_60632
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 46.002 249.792 46.03 ;
      END
   END n_60632

   PIN n_61085
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 32.882 249.792 32.91 ;
      END
   END n_61085

   PIN n_61149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.866 249.792 18.894 ;
      END
   END n_61149

   PIN n_61187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 15.218 249.792 15.246 ;
      END
   END n_61187

   PIN n_61461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.274 117.597 220.302 117.76 ;
      END
   END n_61461

   PIN n_61579
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.058 249.792 11.086 ;
      END
   END n_61579

   PIN n_61580
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.802 249.792 18.83 ;
      END
   END n_61580

   PIN n_61592
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 92.21 249.792 92.238 ;
      END
   END n_61592

   PIN n_61601
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 49.714 249.792 49.742 ;
      END
   END n_61601

   PIN n_61705
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.394 117.597 97.422 117.76 ;
      END
   END n_61705

   PIN n_61723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.25 0.0 51.278 0.163 ;
      END
   END n_61723

   PIN n_61755
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 102.898 0.0 102.926 0.163 ;
      END
   END n_61755

   PIN n_61873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 103.922 249.792 103.95 ;
      END
   END n_61873

   PIN n_61878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.082 117.597 228.11 117.76 ;
      END
   END n_61878

   PIN n_61893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.434 117.597 216.462 117.76 ;
      END
   END n_61893

   PIN n_61956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 8.306 249.792 8.334 ;
      END
   END n_61956

   PIN n_62290
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 60.978 249.792 61.006 ;
      END
   END n_62290

   PIN n_62406
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 65.138 249.792 65.166 ;
      END
   END n_62406

   PIN n_62437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.21 117.597 220.238 117.76 ;
      END
   END n_62437

   PIN n_62460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.594 117.597 212.622 117.76 ;
      END
   END n_62460

   PIN n_62694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 204.85 117.597 204.878 117.76 ;
      END
   END n_62694

   PIN n_62695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 212.722 117.597 212.75 117.76 ;
      END
   END n_62695

   PIN n_63124
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 18.162 249.792 18.19 ;
      END
   END n_63124

   PIN n_63132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 49.394 249.792 49.422 ;
      END
   END n_63132

   PIN n_63155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.458 0.0 89.486 0.163 ;
      END
   END n_63155

   PIN n_63260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 174.258 117.597 174.286 117.76 ;
      END
   END n_63260

   PIN n_63263
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.074 117.597 137.102 117.76 ;
      END
   END n_63263

   PIN n_63360
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.554 0.0 181.582 0.163 ;
      END
   END n_63360

   PIN n_63423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 27.25 249.792 27.278 ;
      END
   END n_63423

   PIN n_63445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 70.514 249.792 70.542 ;
      END
   END n_63445

   PIN n_63901
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.146 117.597 220.174 117.76 ;
      END
   END n_63901

   PIN n_64318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.106 117.597 149.134 117.76 ;
      END
   END n_64318

   PIN n_64366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 11.122 249.792 11.15 ;
      END
   END n_64366

   PIN n_64478
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.962 249.792 62.99 ;
      END
   END n_64478

   PIN n_64560
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.69 117.597 224.718 117.76 ;
      END
   END n_64560

   PIN n_64768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.106 249.792 77.134 ;
      END
   END n_64768

   PIN n_64772
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 80.882 249.792 80.91 ;
      END
   END n_64772

   PIN n_64912
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.002 117.597 150.03 117.76 ;
      END
   END n_64912

   PIN n_65026
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.562 117.597 216.59 117.76 ;
      END
   END n_65026

   PIN n_65319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.602 0.0 87.63 0.163 ;
      END
   END n_65319

   PIN n_65354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.026 117.597 143.054 117.76 ;
      END
   END n_65354

   PIN n_65426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.458 117.597 97.486 117.76 ;
      END
   END n_65426

   PIN n_65480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.794 249.792 47.822 ;
      END
   END n_65480

   PIN n_65483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 54.898 249.792 54.926 ;
      END
   END n_65483

   PIN n_65893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.234 249.792 77.262 ;
      END
   END n_65893

   PIN n_65894
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 77.042 249.792 77.07 ;
      END
   END n_65894

   PIN n_66724
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.53 117.597 212.558 117.76 ;
      END
   END n_66724

   PIN n_66751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.746 249.792 77.774 ;
      END
   END n_66751

   PIN n_66842
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.786 249.792 84.814 ;
      END
   END n_66842

   PIN n_66843
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 84.722 249.792 84.75 ;
      END
   END n_66843

   PIN n_66867
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.042 117.597 149.07 117.76 ;
      END
   END n_66867

   PIN n_67068
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.81 0.0 85.838 0.163 ;
      END
   END n_67068

   PIN n_67215
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 47.73 249.792 47.758 ;
      END
   END n_67215

   PIN n_70345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 91.762 249.792 91.79 ;
      END
   END n_70345

   PIN n_70642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.41 117.597 239.438 117.76 ;
      END
   END n_70642

   PIN n_71222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.442 249.792 99.47 ;
      END
   END n_71222

   PIN n_71449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.162 0.0 98.19 0.163 ;
      END
   END n_71449

   PIN n_71795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.874 0.0 157.902 0.163 ;
      END
   END n_71795

   PIN n_77679
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.41 0.0 143.438 0.163 ;
      END
   END n_77679

   PIN n_77842
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 84.722 0.0 84.75 0.163 ;
      END
   END n_77842

   PIN n_80858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 114.162 249.792 114.19 ;
      END
   END n_80858

   PIN n_81895
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 77.682 249.792 77.71 ;
      END
   END n_81895

   PIN n_82145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.874 117.597 181.902 117.76 ;
      END
   END n_82145

   PIN n_82355
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 88.114 249.792 88.142 ;
      END
   END n_82355

   PIN n_82437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 239.538 117.597 239.566 117.76 ;
      END
   END n_82437

   PIN n_8249
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.058 0.0 51.086 0.163 ;
      END
   END n_8249

   PIN n_82916
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 62.514 249.792 62.542 ;
      END
   END n_82916

   PIN n_83187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 95.858 249.792 95.886 ;
      END
   END n_83187

   PIN n_83203
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.762 249.792 99.79 ;
      END
   END n_83203

   PIN n_84332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 115.122 249.792 115.15 ;
      END
   END n_84332

   PIN n_85306
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 249.629 95.986 249.792 96.014 ;
      END
   END n_85306

   PIN n_85307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 99.634 249.792 99.662 ;
      END
   END n_85307

   PIN n_85541
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 177.97 0.0 177.998 0.163 ;
      END
   END n_85541

   PIN n_86195
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 72.626 249.792 72.654 ;
      END
   END n_86195

   PIN n_87554
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.81 117.597 181.838 117.76 ;
      END
   END n_87554

   PIN n_87555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.746 117.597 181.774 117.76 ;
      END
   END n_87555

   PIN n_88558
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 249.629 95.794 249.792 95.822 ;
      END
   END n_88558

   PIN n_95316
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 248.562 117.597 248.59 117.76 ;
      END
   END n_95316

   PIN n_95932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 32.242 0.0 32.27 0.163 ;
      END
   END n_95932

   PIN n_96299
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.098 117.597 186.126 117.76 ;
      END
   END n_96299

   PIN n_96642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.754 0.0 40.782 0.163 ;
      END
   END n_96642

   PIN n_97723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.218 0.0 151.246 0.163 ;
      END
   END n_97723

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER V1 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 249.792 117.76 ;
      LAYER M1 ;
         RECT 0.0 0.0 249.792 117.76 ;
   END
END h2_mgc_matrix_mult_b

MACRO h1_mgc_matrix_mult_b
   CLASS BLOCK ;
   FOREIGN h1 ;
   ORIGIN 0 0 ;
   SIZE 257.902 BY 159.362 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN15738_FE_OFN11549_n_142793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.778 159.198 113.806 159.362 ;
      END
   END FE_OCPN15738_FE_OFN11549_n_142793

   PIN FE_OFN10667_a_5_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 126.706 257.902 126.734 ;
      END
   END FE_OFN10667_a_5_6_4

   PIN FE_OFN10748_a_4_4_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 80.562 257.902 80.59 ;
      END
   END FE_OFN10748_a_4_4_4

   PIN FE_OFN10792_a_4_0_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 88.37 257.902 88.398 ;
      END
   END FE_OFN10792_a_4_0_5

   PIN FE_OFN10799_a_3_8_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 134.194 257.902 134.222 ;
      END
   END FE_OFN10799_a_3_8_7

   PIN FE_OFN10820_a_3_6_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 104.562 257.902 104.59 ;
      END
   END FE_OFN10820_a_3_6_7

   PIN FE_OFN10830_a_3_4_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 85.362 257.902 85.39 ;
      END
   END FE_OFN10830_a_3_4_5

   PIN FE_OFN10834_a_3_4_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 92.21 257.902 92.238 ;
      END
   END FE_OFN10834_a_3_4_0

   PIN FE_OFN10851_a_2_8_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 92.786 257.902 92.814 ;
      END
   END FE_OFN10851_a_2_8_4

   PIN FE_OFN10859_a_2_8_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 123.698 257.902 123.726 ;
      END
   END FE_OFN10859_a_2_8_1

   PIN FE_OFN10872_a_2_6_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 80.626 257.902 80.654 ;
      END
   END FE_OFN10872_a_2_6_7

   PIN FE_OFN10879_a_2_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 92.274 257.902 92.302 ;
      END
   END FE_OFN10879_a_2_6_4

   PIN FE_OFN10888_a_2_4_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 114.354 257.902 114.382 ;
      END
   END FE_OFN10888_a_2_4_7

   PIN FE_OFN10898_a_2_4_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 214.514 0.0 214.542 0.163 ;
      END
   END FE_OFN10898_a_2_4_1

   PIN FE_OFN10902_a_2_4_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 84.338 257.902 84.366 ;
      END
   END FE_OFN10902_a_2_4_0

   PIN FE_OFN10931_a_1_4_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 92.85 257.902 92.878 ;
      END
   END FE_OFN10931_a_1_4_0

   PIN FE_OFN10982_a_0_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 143.666 257.902 143.694 ;
      END
   END FE_OFN10982_a_0_6_4

   PIN FE_OFN10987_a_0_6_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 95.858 257.902 95.886 ;
      END
   END FE_OFN10987_a_0_6_1

   PIN FE_OFN10999_a_0_4_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.426 257.902 85.454 ;
      END
   END FE_OFN10999_a_0_4_7

   PIN FE_OFN11007_a_0_4_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 80.754 257.902 80.782 ;
      END
   END FE_OFN11007_a_0_4_0

   PIN FE_OFN12751_n_142961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.162 159.198 90.19 159.362 ;
      END
   END FE_OFN12751_n_142961

   PIN FE_OFN12753_n_142961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.122 159.198 123.15 159.362 ;
      END
   END FE_OFN12753_n_142961

   PIN FE_OFN14480_n_112183
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.546 159.198 154.574 159.362 ;
      END
   END FE_OFN14480_n_112183

   PIN FE_OFN14491_n_112182
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.074 159.198 121.102 159.362 ;
      END
   END FE_OFN14491_n_112182

   PIN FE_OFN14493_n_112182
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.698 159.198 147.726 159.362 ;
      END
   END FE_OFN14493_n_112182

   PIN FE_OFN14699_a_9_6_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 123.762 257.902 123.79 ;
      END
   END FE_OFN14699_a_9_6_7

   PIN FE_OFN14911_n_142849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.842 159.198 97.87 159.362 ;
      END
   END FE_OFN14911_n_142849

   PIN FE_OFN15367_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.586 159.198 201.614 159.362 ;
      END
   END FE_OFN15367_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_13_

   PIN FE_OFN15376_n_21671
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 157.426 257.902 157.454 ;
      END
   END FE_OFN15376_n_21671

   PIN FE_OFN15983_n_36821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.394 159.198 105.422 159.362 ;
      END
   END FE_OFN15983_n_36821

   PIN FE_OFN16026_a_0_6_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 73.01 257.902 73.038 ;
      END
   END FE_OFN16026_a_0_6_1

   PIN FE_OFN16151_a_2_4_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 75.89 257.902 75.918 ;
      END
   END FE_OFN16151_a_2_4_5

   PIN FE_OFN16443_a_7_4_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.49 257.902 85.518 ;
      END
   END FE_OFN16443_a_7_4_5

   PIN FE_OFN16476_a_2_6_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 217.01 0.0 217.038 0.163 ;
      END
   END FE_OFN16476_a_2_6_1

   PIN FE_OFN17481_n_126984
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.682 0.0 101.71 0.163 ;
      END
   END FE_OFN17481_n_126984

   PIN FE_OFN17555_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.818 159.198 120.846 159.362 ;
      END
   END FE_OFN17555_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_

   PIN FE_OFN18498_n_22234
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.914 159.198 212.942 159.362 ;
      END
   END FE_OFN18498_n_22234

   PIN FE_OFN18638_a_7_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 88.306 257.902 88.334 ;
      END
   END FE_OFN18638_a_7_6_4

   PIN FE_OFN18656_a_3_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 88.37 257.902 88.398 ;
      END
   END FE_OFN18656_a_3_6_4

   PIN FE_OFN18679_a_1_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 134.258 257.902 134.286 ;
      END
   END FE_OFN18679_a_1_6_4

   PIN FE_OFN19318_a_8_8_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 143.73 257.902 143.758 ;
      END
   END FE_OFN19318_a_8_8_4

   PIN FE_OFN19321_a_4_6_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 92.914 257.902 92.942 ;
      END
   END FE_OFN19321_a_4_6_4

   PIN FE_OFN437_n_21145
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 157.49 257.902 157.518 ;
      END
   END FE_OFN437_n_21145

   PIN FE_OFN4661_n_142849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.93 159.198 74.958 159.362 ;
      END
   END FE_OFN4661_n_142849

   PIN FE_OFN4678_n_112357
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.97 159.198 89.998 159.362 ;
      END
   END FE_OFN4678_n_112357

   PIN FE_OFN4703_n_143619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.754 159.198 120.782 159.362 ;
      END
   END FE_OFN4703_n_143619

   PIN FE_OFN4840_n_140222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 143.986 159.198 144.014 159.362 ;
      END
   END FE_OFN4840_n_140222

   PIN FE_OFN4981_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 232.242 159.198 232.27 159.362 ;
      END
   END FE_OFN4981_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_11_

   PIN FE_OFN4983_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 236.146 159.198 236.174 159.362 ;
      END
   END FE_OFN4983_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_10_

   PIN FE_OFN5000_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 245.17 159.198 245.198 159.362 ;
      END
   END FE_OFN5000_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_11_

   PIN FE_OFN636_n_11194
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 92.018 257.902 92.046 ;
      END
   END FE_OFN636_n_11194

   PIN FE_OFN638_n_8336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 7.858 257.902 7.886 ;
      END
   END FE_OFN638_n_8336

   PIN FE_OFN651_n_7003
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 213.106 0.0 213.134 0.163 ;
      END
   END FE_OFN651_n_7003

   PIN FE_OFN741_n_22817
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.01 0.0 121.038 0.163 ;
      END
   END FE_OFN741_n_22817

   PIN FE_OFN8951_n_6635
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.642 159.198 150.67 159.362 ;
      END
   END FE_OFN8951_n_6635

   PIN FE_OFN9215_delay_add_ln34_unr2_unr8_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 17.458 257.902 17.486 ;
      END
   END FE_OFN9215_delay_add_ln34_unr2_unr8_stage2_stallmux_q_13_

   PIN FE_OFN9217_delay_add_ln34_unr2_unr8_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 75.954 257.902 75.982 ;
      END
   END FE_OFN9217_delay_add_ln34_unr2_unr8_stage2_stallmux_q_12_

   PIN FE_OFN9884_b_4_8_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.146 159.198 4.174 159.362 ;
      END
   END FE_OFN9884_b_4_8_1

   PIN FE_OFN9902_b_4_7_9
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.778 159.198 97.806 159.362 ;
      END
   END FE_OFN9902_b_4_7_9

   PIN delay_add_ln34_unr2_unr1_stage2_stallmux_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 7.922 257.902 7.95 ;
      END
   END delay_add_ln34_unr2_unr1_stage2_stallmux_q_10_

   PIN delay_add_ln34_unr2_unr1_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 17.522 257.902 17.55 ;
      END
   END delay_add_ln34_unr2_unr1_stage2_stallmux_q_7_

   PIN delay_add_ln34_unr2_unr2_stage2_stallmux_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 145.842 257.902 145.87 ;
      END
   END delay_add_ln34_unr2_unr2_stage2_stallmux_q_1_

   PIN delay_add_ln34_unr2_unr2_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 37.426 257.902 37.454 ;
      END
   END delay_add_ln34_unr2_unr2_stage2_stallmux_q_2_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 17.586 257.902 17.614 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_12_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 206.706 0.0 206.734 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_14_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.106 0.0 117.134 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_7_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.042 0.0 117.07 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr3_unr7_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.618 159.198 101.646 159.362 ;
      END
   END delay_mul_ln34_unr3_unr7_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.578 159.198 166.606 159.362 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr4_unr7_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.322 0.0 182.35 0.163 ;
      END
   END delay_mul_ln34_unr4_unr7_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr4_unr9_stage2_stallmux_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 107.57 257.902 107.598 ;
      END
   END delay_mul_ln34_unr4_unr9_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.922 159.198 239.95 159.362 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 232.306 159.198 232.334 159.362 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_13_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.786 159.198 220.814 159.362 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_14_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 236.21 159.198 236.238 159.362 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.45 159.198 182.478 159.362 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.442 159.198 155.47 159.362 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_9_

   PIN mul_4646_72_n_150
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.682 159.198 101.71 159.362 ;
      END
   END mul_4646_72_n_150

   PIN mul_4646_72_n_251
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.01 159.198 121.038 159.362 ;
      END
   END mul_4646_72_n_251

   PIN mul_4646_72_n_58
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.522 0.0 105.55 0.163 ;
      END
   END mul_4646_72_n_58

   PIN mul_4646_72_n_59
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.33 0.0 113.358 0.163 ;
      END
   END mul_4646_72_n_59

   PIN mul_4646_72_n_75
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.122 0.0 115.15 0.163 ;
      END
   END mul_4646_72_n_75

   PIN mul_4646_72_n_756
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.514 0.0 134.542 0.163 ;
      END
   END mul_4646_72_n_756

   PIN mul_4650_72_n_212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.594 159.198 132.622 159.362 ;
      END
   END mul_4650_72_n_212

   PIN mul_4650_72_n_213
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.402 159.198 132.43 159.362 ;
      END
   END mul_4650_72_n_213

   PIN mul_4650_72_n_214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 141.298 159.198 141.326 159.362 ;
      END
   END mul_4650_72_n_214

   PIN mul_4650_72_n_217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.21 0.0 44.238 0.163 ;
      END
   END mul_4650_72_n_217

   PIN mul_4650_72_n_239
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.802 159.198 74.83 159.362 ;
      END
   END mul_4650_72_n_239

   PIN mul_4650_72_n_252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.146 159.198 36.174 159.362 ;
      END
   END mul_4650_72_n_252

   PIN mul_4650_72_n_285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 67.058 159.198 67.086 159.362 ;
      END
   END mul_4650_72_n_285

   PIN mul_4650_72_n_287
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.834 159.198 70.862 159.362 ;
      END
   END mul_4650_72_n_287

   PIN mul_4650_72_n_289
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.442 159.198 59.47 159.362 ;
      END
   END mul_4650_72_n_289

   PIN mul_4650_72_n_292
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.37 159.198 40.398 159.362 ;
      END
   END mul_4650_72_n_292

   PIN mul_4650_72_n_311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 86.77 159.198 86.798 159.362 ;
      END
   END mul_4650_72_n_311

   PIN mul_4650_72_n_313
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.482 159.198 82.51 159.362 ;
      END
   END mul_4650_72_n_313

   PIN mul_4650_72_n_55
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.954 0.0 51.982 0.163 ;
      END
   END mul_4650_72_n_55

   PIN mul_4650_72_n_73
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.674 0.0 106.702 0.163 ;
      END
   END mul_4650_72_n_73

   PIN mul_4650_72_n_777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.018 0.0 52.046 0.163 ;
      END
   END mul_4650_72_n_777

   PIN mul_4650_72_n_78
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.466 159.198 132.494 159.362 ;
      END
   END mul_4650_72_n_78

   PIN mul_4650_72_n_848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.17 0.0 53.198 0.163 ;
      END
   END mul_4650_72_n_848

   PIN n_111907
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.53 159.198 132.558 159.362 ;
      END
   END n_111907

   PIN n_112284
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.402 159.198 36.43 159.362 ;
      END
   END n_112284

   PIN n_112720
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 132.402 159.198 132.43 159.362 ;
      END
   END n_112720

   PIN n_113639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.122 159.198 51.15 159.362 ;
      END
   END n_113639

   PIN n_113790
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.546 159.198 82.574 159.362 ;
      END
   END n_113790

   PIN n_114086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.946 159.198 120.974 159.362 ;
      END
   END n_114086

   PIN n_114387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.13 0.0 94.158 0.163 ;
      END
   END n_114387

   PIN n_114392
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.058 159.198 51.086 159.362 ;
      END
   END n_114392

   PIN n_114607
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.834 0.0 94.862 0.163 ;
      END
   END n_114607

   PIN n_114644
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.37 159.198 120.398 159.362 ;
      END
   END n_114644

   PIN n_114654
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.346 159.198 63.374 159.362 ;
      END
   END n_114654

   PIN n_115067
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.706 0.0 78.734 0.163 ;
      END
   END n_115067

   PIN n_115075
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.73 0.0 55.758 0.163 ;
      END
   END n_115075

   PIN n_115173
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.666 0.0 55.694 0.163 ;
      END
   END n_115173

   PIN n_115193
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.354 159.198 106.382 159.362 ;
      END
   END n_115193

   PIN n_115538
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 118.706 159.198 118.734 159.362 ;
      END
   END n_115538

   PIN n_115592
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.41 159.198 63.438 159.362 ;
      END
   END n_115592

   PIN n_115601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.81 159.198 93.838 159.362 ;
      END
   END n_115601

   PIN n_115610
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.682 159.198 101.71 159.362 ;
      END
   END n_115610

   PIN n_115697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.65 159.198 105.678 159.362 ;
      END
   END n_115697

   PIN n_115863
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.706 159.198 30.734 159.362 ;
      END
   END n_115863

   PIN n_115878
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.482 159.198 58.51 159.362 ;
      END
   END n_115878

   PIN n_115897
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.482 159.198 34.51 159.362 ;
      END
   END n_115897

   PIN n_116017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.522 159.198 105.55 159.362 ;
      END
   END n_116017

   PIN n_116364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.426 159.198 101.454 159.362 ;
      END
   END n_116364

   PIN n_116388
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.41 159.198 63.438 159.362 ;
      END
   END n_116388

   PIN n_116530
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.746 159.198 101.774 159.362 ;
      END
   END n_116530

   PIN n_116580
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.066 159.198 94.094 159.362 ;
      END
   END n_116580

   PIN n_116853
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.362 159.198 109.39 159.362 ;
      END
   END n_116853

   PIN n_116869
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.258 159.198 94.286 159.362 ;
      END
   END n_116869

   PIN n_117308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.146 0.0 44.174 0.163 ;
      END
   END n_117308

   PIN n_117932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.834 159.198 46.862 159.362 ;
      END
   END n_117932

   PIN n_118446
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.874 159.198 117.902 159.362 ;
      END
   END n_118446

   PIN n_118851
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.29 159.198 50.318 159.362 ;
      END
   END n_118851

   PIN n_118961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 96.754 159.198 96.782 159.362 ;
      END
   END n_118961

   PIN n_119042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.858 159.198 103.886 159.362 ;
      END
   END n_119042

   PIN n_119323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 98.098 159.198 98.126 159.362 ;
      END
   END n_119323

   PIN n_119415
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.506 159.198 107.534 159.362 ;
      END
   END n_119415

   PIN n_119457
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.186 159.198 67.214 159.362 ;
      END
   END n_119457

   PIN n_120207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.33 159.198 113.358 159.362 ;
      END
   END n_120207

   PIN n_120352
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.77 0.0 78.798 0.163 ;
      END
   END n_120352

   PIN n_120375
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.498 159.198 120.526 159.362 ;
      END
   END n_120375

   PIN n_120599
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.426 0.0 109.454 0.163 ;
      END
   END n_120599

   PIN n_120600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.81 0.0 101.838 0.163 ;
      END
   END n_120600

   PIN n_121035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.746 159.198 117.774 159.362 ;
      END
   END n_121035

   PIN n_121273
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.21 0.0 44.238 0.163 ;
      END
   END n_121273

   PIN n_121548
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.33 159.198 17.358 159.362 ;
      END
   END n_121548

   PIN n_121555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 98.034 159.198 98.062 159.362 ;
      END
   END n_121555

   PIN n_121639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.722 159.198 124.75 159.362 ;
      END
   END n_121639

   PIN n_121887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.794 0.0 63.822 0.163 ;
      END
   END n_121887

   PIN n_121951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.45 0.0 86.478 0.163 ;
      END
   END n_121951

   PIN n_122050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.514 0.0 86.542 0.163 ;
      END
   END n_122050

   PIN n_122090
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.666 159.198 55.694 159.362 ;
      END
   END n_122090

   PIN n_122254
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.506 0.0 59.534 0.163 ;
      END
   END n_122254

   PIN n_122427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 88.498 257.902 88.526 ;
      END
   END n_122427

   PIN n_124381
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 99.89 257.902 99.918 ;
      END
   END n_124381

   PIN n_124384
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.554 257.902 85.582 ;
      END
   END n_124384

   PIN n_124473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.922 0.0 47.95 0.163 ;
      END
   END n_124473

   PIN n_124480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.178 159.198 24.206 159.362 ;
      END
   END n_124480

   PIN n_124768
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.674 159.198 138.702 159.362 ;
      END
   END n_124768

   PIN n_124884
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.01 159.198 129.038 159.362 ;
      END
   END n_124884

   PIN n_124890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.882 159.198 120.91 159.362 ;
      END
   END n_124890

   PIN n_124892
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.906 0.0 97.934 0.163 ;
      END
   END n_124892

   PIN n_125201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 92.338 257.902 92.366 ;
      END
   END n_125201

   PIN n_125438
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.266 0.0 113.294 0.163 ;
      END
   END n_125438

   PIN n_125484
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.714 0.0 89.742 0.163 ;
      END
   END n_125484

   PIN n_126152
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 92.082 257.902 92.11 ;
      END
   END n_126152

   PIN n_126230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 88.434 257.902 88.462 ;
      END
   END n_126230

   PIN n_126465
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.594 0.0 124.622 0.163 ;
      END
   END n_126465

   PIN n_126950
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.69 159.198 32.718 159.362 ;
      END
   END n_126950

   PIN n_127100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.074 0.0 65.102 0.163 ;
      END
   END n_127100

   PIN n_127101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.01 0.0 65.038 0.163 ;
      END
   END n_127101

   PIN n_127102
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.282 0.0 63.31 0.163 ;
      END
   END n_127102

   PIN n_127132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.258 159.198 126.286 159.362 ;
      END
   END n_127132

   PIN n_127133
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.194 159.198 126.222 159.362 ;
      END
   END n_127133

   PIN n_127136
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.97 0.0 97.998 0.163 ;
      END
   END n_127136

   PIN n_127563
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.69 0.0 128.718 0.163 ;
      END
   END n_127563

   PIN n_128225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.666 0.0 55.694 0.163 ;
      END
   END n_128225

   PIN n_129278
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.986 0.0 48.014 0.163 ;
      END
   END n_129278

   PIN n_130041
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.178 0.0 48.206 0.163 ;
      END
   END n_130041

   PIN n_130821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.642 0.0 22.67 0.163 ;
      END
   END n_130821

   PIN n_131531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.57 0.0 59.598 0.163 ;
      END
   END n_131531

   PIN n_133774
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.89 0.0 51.918 0.163 ;
      END
   END n_133774

   PIN n_13498
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.522 159.198 161.55 159.362 ;
      END
   END n_13498

   PIN n_137441
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.442 0.0 139.47 0.163 ;
      END
   END n_137441

   PIN n_142793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 132.466 159.198 132.494 159.362 ;
      END
   END n_142793

   PIN n_142961
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 103.538 257.902 103.566 ;
      END
   END n_142961

   PIN n_143003
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.538 159.198 63.566 159.362 ;
      END
   END n_143003

   PIN n_14932
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 194.674 159.198 194.702 159.362 ;
      END
   END n_14932

   PIN n_14933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 188.914 159.198 188.942 159.362 ;
      END
   END n_14933

   PIN n_14966
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 190.258 159.198 190.286 159.362 ;
      END
   END n_14966

   PIN n_16625
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.618 257.902 85.646 ;
      END
   END n_16625

   PIN n_16626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.81 257.902 85.838 ;
      END
   END n_16626

   PIN n_17619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 111.346 257.902 111.374 ;
      END
   END n_17619

   PIN n_19300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 151.73 159.198 151.758 159.362 ;
      END
   END n_19300

   PIN n_19852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.21 159.198 196.238 159.362 ;
      END
   END n_19852

   PIN n_19853
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.226 159.198 186.254 159.362 ;
      END
   END n_19853

   PIN n_20189
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.234 0.0 229.262 0.163 ;
      END
   END n_20189

   PIN n_20626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.962 159.198 166.99 159.362 ;
      END
   END n_20626

   PIN n_21390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 85.298 257.902 85.326 ;
      END
   END n_21390

   PIN n_21391
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.682 257.902 85.71 ;
      END
   END n_21391

   PIN n_21448
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.274 159.198 164.302 159.362 ;
      END
   END n_21448

   PIN n_21461
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 174.706 0.0 174.734 0.163 ;
      END
   END n_21461

   PIN n_21505
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.362 159.198 205.39 159.362 ;
      END
   END n_21505

   PIN n_21517
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 138.226 257.902 138.254 ;
      END
   END n_21517

   PIN n_21590
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 179.058 159.198 179.086 159.362 ;
      END
   END n_21590

   PIN n_21591
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 167.026 159.198 167.054 159.362 ;
      END
   END n_21591

   PIN n_21678
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 158.514 159.198 158.542 159.362 ;
      END
   END n_21678

   PIN n_21692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 157.362 257.902 157.39 ;
      END
   END n_21692

   PIN n_21696
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.682 159.198 197.71 159.362 ;
      END
   END n_21696

   PIN n_21711
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 76.018 257.902 76.046 ;
      END
   END n_21711

   PIN n_21955
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.554 0.0 109.582 0.163 ;
      END
   END n_21955

   PIN n_21973
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 209.33 159.198 209.358 159.362 ;
      END
   END n_21973

   PIN n_21974
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 213.042 159.198 213.07 159.362 ;
      END
   END n_21974

   PIN n_21990
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.154 0.0 231.182 0.163 ;
      END
   END n_21990

   PIN n_22100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.49 0.0 109.518 0.163 ;
      END
   END n_22100

   PIN n_22130
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.298 159.198 205.326 159.362 ;
      END
   END n_22130

   PIN n_22131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.426 159.198 205.454 159.362 ;
      END
   END n_22131

   PIN n_22132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.826 159.198 195.854 159.362 ;
      END
   END n_22132

   PIN n_22135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 209.33 159.198 209.358 159.362 ;
      END
   END n_22135

   PIN n_22222
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 243.762 159.198 243.79 159.362 ;
      END
   END n_22222

   PIN n_22223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 159.346 159.198 159.374 159.362 ;
      END
   END n_22223

   PIN n_22241
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 69.042 257.902 69.07 ;
      END
   END n_22241

   PIN n_22502
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.17 0.0 117.198 0.163 ;
      END
   END n_22502

   PIN n_22542
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 45.938 257.902 45.966 ;
      END
   END n_22542

   PIN n_23096
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 138.29 257.902 138.318 ;
      END
   END n_23096

   PIN n_23324
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 119.026 257.902 119.054 ;
      END
   END n_23324

   PIN n_23325
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 17.65 257.902 17.678 ;
      END
   END n_23325

   PIN n_23968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.49 159.198 205.518 159.362 ;
      END
   END n_23968

   PIN n_23969
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.474 159.198 199.502 159.362 ;
      END
   END n_23969

   PIN n_23973
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.65 159.198 201.678 159.362 ;
      END
   END n_23973

   PIN n_24209
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.506 159.198 155.534 159.362 ;
      END
   END n_24209

   PIN n_24210
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.602 159.198 151.63 159.362 ;
      END
   END n_24210

   PIN n_24293
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 119.09 257.902 119.118 ;
      END
   END n_24293

   PIN n_24393
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 157.554 257.902 157.582 ;
      END
   END n_24393

   PIN n_24834
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.058 159.198 155.086 159.362 ;
      END
   END n_24834

   PIN n_24836
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.61 159.198 154.638 159.362 ;
      END
   END n_24836

   PIN n_24845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.034 159.198 146.062 159.362 ;
      END
   END n_24845

   PIN n_24847
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.906 159.198 145.934 159.362 ;
      END
   END n_24847

   PIN n_24890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 209.202 159.198 209.23 159.362 ;
      END
   END n_24890

   PIN n_24892
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 209.266 159.198 209.294 159.362 ;
      END
   END n_24892

   PIN n_24997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 141.874 257.902 141.902 ;
      END
   END n_24997

   PIN n_25050
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 134.386 257.902 134.414 ;
      END
   END n_25050

   PIN n_25074
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 155.57 159.198 155.598 159.362 ;
      END
   END n_25074

   PIN n_25101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 209.394 159.198 209.422 159.362 ;
      END
   END n_25101

   PIN n_25132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 114.994 257.902 115.022 ;
      END
   END n_25132

   PIN n_25257
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 149.234 159.198 149.262 159.362 ;
      END
   END n_25257

   PIN n_25529
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.666 159.198 151.694 159.362 ;
      END
   END n_25529

   PIN n_25531
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 151.666 159.198 151.694 159.362 ;
      END
   END n_25531

   PIN n_25624
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 111.41 257.902 111.438 ;
      END
   END n_25624

   PIN n_26550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 197.81 159.198 197.838 159.362 ;
      END
   END n_26550

   PIN n_26818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.746 159.198 197.774 159.362 ;
      END
   END n_26818

   PIN n_27649
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.026 159.198 231.054 159.362 ;
      END
   END n_27649

   PIN n_27650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 232.37 159.198 232.398 159.362 ;
      END
   END n_27650

   PIN n_27752
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 217.01 159.198 217.038 159.362 ;
      END
   END n_27752

   PIN n_2800
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.05 0.0 48.078 0.163 ;
      END
   END n_2800

   PIN n_28028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.626 159.198 224.654 159.362 ;
      END
   END n_28028

   PIN n_28030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.53 159.198 228.558 159.362 ;
      END
   END n_28030

   PIN n_28637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.85 159.198 220.878 159.362 ;
      END
   END n_28637

   PIN n_28704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 174.77 0.0 174.798 0.163 ;
      END
   END n_28704

   PIN n_28825
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 251.698 159.198 251.726 159.362 ;
      END
   END n_28825

   PIN n_29574
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 145.906 257.902 145.934 ;
      END
   END n_29574

   PIN n_29646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 143.794 257.902 143.822 ;
      END
   END n_29646

   PIN n_32056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.258 159.198 78.286 159.362 ;
      END
   END n_32056

   PIN n_32073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.05 159.198 88.078 159.362 ;
      END
   END n_32073

   PIN n_32468
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.33 159.198 113.358 159.362 ;
      END
   END n_32468

   PIN n_32697
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.802 159.198 170.83 159.362 ;
      END
   END n_32697

   PIN n_32704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.434 159.198 40.462 159.362 ;
      END
   END n_32704

   PIN n_32867
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.866 159.198 170.894 159.362 ;
      END
   END n_32867

   PIN n_33365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.93 159.198 170.958 159.362 ;
      END
   END n_33365

   PIN n_33776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.226 159.198 130.254 159.362 ;
      END
   END n_33776

   PIN n_34364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.474 159.198 63.502 159.362 ;
      END
   END n_34364

   PIN n_34374
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.602 159.198 55.63 159.362 ;
      END
   END n_34374

   PIN n_34614
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 104.37 159.198 104.398 159.362 ;
      END
   END n_34614

   PIN n_34686
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 129.97 159.198 129.998 159.362 ;
      END
   END n_34686

   PIN n_35435
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.21 159.198 44.238 159.362 ;
      END
   END n_35435

   PIN n_35467
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.93 159.198 106.958 159.362 ;
      END
   END n_35467

   PIN n_36948
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.434 159.198 72.462 159.362 ;
      END
   END n_36948

   PIN n_37020
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.314 159.198 67.342 159.362 ;
      END
   END n_37020

   PIN n_37253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.866 159.198 74.894 159.362 ;
      END
   END n_37253

   PIN n_37497
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.522 159.198 25.55 159.362 ;
      END
   END n_37497

   PIN n_37498
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.89 159.198 19.918 159.362 ;
      END
   END n_37498

   PIN n_37637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.322 159.198 110.35 159.362 ;
      END
   END n_37637

   PIN n_38077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.074 0.0 113.102 0.163 ;
      END
   END n_38077

   PIN n_39307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.746 0.0 101.774 0.163 ;
      END
   END n_39307

   PIN n_39821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 134.322 257.902 134.35 ;
      END
   END n_39821

   PIN n_39967
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 46.962 257.902 46.99 ;
      END
   END n_39967

   PIN n_40268
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 80.562 257.902 80.59 ;
      END
   END n_40268

   PIN n_40473
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 76.082 257.902 76.11 ;
      END
   END n_40473

   PIN n_40638
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 80.626 257.902 80.654 ;
      END
   END n_40638

   PIN n_40714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 88.178 257.902 88.206 ;
      END
   END n_40714

   PIN n_41448
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.858 159.198 143.886 159.362 ;
      END
   END n_41448

   PIN n_44877
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.93 159.198 74.958 159.362 ;
      END
   END n_44877

   PIN n_47745
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.186 159.198 91.214 159.362 ;
      END
   END n_47745

   PIN n_47887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.546 159.198 82.574 159.362 ;
      END
   END n_47887

   PIN n_48179
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.034 159.198 74.062 159.362 ;
      END
   END n_48179

   PIN n_54122
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.898 159.198 70.926 159.362 ;
      END
   END n_54122

   PIN n_54294
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.25 159.198 67.278 159.362 ;
      END
   END n_54294

   PIN n_5456
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.93 0.0 106.958 0.163 ;
      END
   END n_5456

   PIN n_5457
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.378 0.0 107.406 0.163 ;
      END
   END n_5457

   PIN n_57601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.562 159.198 72.59 159.362 ;
      END
   END n_57601

   PIN n_59902
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.898 159.198 54.926 159.362 ;
      END
   END n_59902

   PIN n_60533
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.37 159.198 72.398 159.362 ;
      END
   END n_60533

   PIN n_62170
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.61 159.198 74.638 159.362 ;
      END
   END n_62170

   PIN n_6519
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.098 159.198 242.126 159.362 ;
      END
   END n_6519

   PIN n_65559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 219.506 159.198 219.534 159.362 ;
      END
   END n_65559

   PIN n_7333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 178.61 0.0 178.638 0.163 ;
      END
   END n_7333

   PIN n_8253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 53.746 257.902 53.774 ;
      END
   END n_8253

   PIN n_9777
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.378 159.198 195.406 159.362 ;
      END
   END n_9777

   PIN FE_OCPN15632_n_40178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 72.946 257.902 72.974 ;
      END
   END FE_OCPN15632_n_40178

   PIN FE_OFN10061_b_4_3_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.418 159.198 74.446 159.362 ;
      END
   END FE_OFN10061_b_4_3_6

   PIN FE_OFN10064_b_4_3_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.898 159.198 110.926 159.362 ;
      END
   END FE_OFN10064_b_4_3_5

   PIN FE_OFN10067_b_4_3_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.306 159.198 88.334 159.362 ;
      END
   END FE_OFN10067_b_4_3_4

   PIN FE_OFN10070_b_4_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 99.826 159.198 99.854 159.362 ;
      END
   END FE_OFN10070_b_4_3_3

   PIN FE_OFN10072_b_4_3_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.474 159.198 111.502 159.362 ;
      END
   END FE_OFN10072_b_4_3_2

   PIN FE_OFN10076_b_4_3_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.026 159.198 95.054 159.362 ;
      END
   END FE_OFN10076_b_4_3_1

   PIN FE_OFN10077_b_4_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.906 159.198 97.934 159.362 ;
      END
   END FE_OFN10077_b_4_3_0

   PIN FE_OFN10078_b_4_3_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.81 159.198 117.838 159.362 ;
      END
   END FE_OFN10078_b_4_3_0

   PIN FE_OFN10180_b_4_0_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.61 159.28 66.638 159.362 ;
      END
   END FE_OFN10180_b_4_0_3

   PIN FE_OFN10188_b_4_0_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.066 159.198 94.094 159.362 ;
      END
   END FE_OFN10188_b_4_0_0

   PIN FE_OFN10818_a_3_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 247.666 159.198 247.694 159.362 ;
      END
   END FE_OFN10818_a_3_6_7

   PIN FE_OFN10857_a_2_8_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 251.57 159.198 251.598 159.362 ;
      END
   END FE_OFN10857_a_2_8_1

   PIN FE_OFN10871_a_2_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.042 159.198 245.07 159.362 ;
      END
   END FE_OFN10871_a_2_6_7

   PIN FE_OFN10986_a_0_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 240.754 159.198 240.782 159.362 ;
      END
   END FE_OFN10986_a_0_6_1

   PIN FE_OFN11519_n_40714
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 95.026 257.902 95.054 ;
      END
   END FE_OFN11519_n_40714

   PIN FE_OFN11549_n_142793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.042 159.198 117.07 159.362 ;
      END
   END FE_OFN11549_n_142793

   PIN FE_OFN1154_n_10378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.666 0.0 151.694 0.163 ;
      END
   END FE_OFN1154_n_10378

   PIN FE_OFN11610_n_39244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.074 159.198 137.102 159.362 ;
      END
   END FE_OFN11610_n_39244

   PIN FE_OFN11880_n_143202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 110.834 159.198 110.862 159.362 ;
      END
   END FE_OFN11880_n_143202

   PIN FE_OFN11883_n_143200
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.866 159.198 74.894 159.362 ;
      END
   END FE_OFN11883_n_143200

   PIN FE_OFN12031_n_143507
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 83.89 159.198 83.918 159.362 ;
      END
   END FE_OFN12031_n_143507

   PIN FE_OFN12057_n_140222
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.674 159.198 82.702 159.362 ;
      END
   END FE_OFN12057_n_140222

   PIN FE_OFN12086_n_143619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.002 159.198 94.03 159.362 ;
      END
   END FE_OFN12086_n_143619

   PIN FE_OFN12427_n_143003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.834 159.198 78.862 159.362 ;
      END
   END FE_OFN12427_n_143003

   PIN FE_OFN12759_n_142961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.258 159.198 110.286 159.362 ;
      END
   END FE_OFN12759_n_142961

   PIN FE_OFN13003_n_39130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.874 159.198 109.902 159.362 ;
      END
   END FE_OFN13003_n_39130

   PIN FE_OFN13192_n_37615
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.482 159.198 82.51 159.362 ;
      END
   END FE_OFN13192_n_37615

   PIN FE_OFN13223_n_143620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.57 159.198 91.598 159.362 ;
      END
   END FE_OFN13223_n_143620

   PIN FE_OFN13288_n_143034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.418 159.198 90.446 159.362 ;
      END
   END FE_OFN13288_n_143034

   PIN FE_OFN13294_n_143033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.306 159.198 120.334 159.362 ;
      END
   END FE_OFN13294_n_143033

   PIN FE_OFN13296_n_143032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.018 159.198 92.046 159.362 ;
      END
   END FE_OFN13296_n_143032

   PIN FE_OFN13353_n_142795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.842 159.198 113.87 159.362 ;
      END
   END FE_OFN13353_n_142795

   PIN FE_OFN13512_n_112357
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.162 159.198 90.19 159.362 ;
      END
   END FE_OFN13512_n_112357

   PIN FE_OFN13586_n_143006
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.738 159.198 74.766 159.362 ;
      END
   END FE_OFN13586_n_143006

   PIN FE_OFN14074_n_142964
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.954 159.198 107.982 159.362 ;
      END
   END FE_OFN14074_n_142964

   PIN FE_OFN14079_n_142963
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.242 159.198 88.27 159.362 ;
      END
   END FE_OFN14079_n_142963

   PIN FE_OFN14083_n_142962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.338 159.198 60.366 159.362 ;
      END
   END FE_OFN14083_n_142962

   PIN FE_OFN14327_n_140207
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.522 159.28 105.55 159.362 ;
      END
   END FE_OFN14327_n_140207

   PIN FE_OFN14360_n_143300
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.698 159.198 51.726 159.362 ;
      END
   END FE_OFN14360_n_143300

   PIN FE_OFN14403_n_142794
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.114 159.28 88.142 159.362 ;
      END
   END FE_OFN14403_n_142794

   PIN FE_OFN14479_n_112183
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.626 159.198 128.654 159.362 ;
      END
   END FE_OFN14479_n_112183

   PIN FE_OFN14487_n_143005
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 102.77 159.198 102.798 159.362 ;
      END
   END FE_OFN14487_n_143005

   PIN FE_OFN14698_a_9_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.962 159.198 246.99 159.362 ;
      END
   END FE_OFN14698_a_9_6_7

   PIN FE_OFN14912_n_142849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.034 159.198 90.062 159.362 ;
      END
   END FE_OFN14912_n_142849

   PIN FE_OFN14984_n_112030
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.81 159.198 101.838 159.362 ;
      END
   END FE_OFN14984_n_112030

   PIN FE_OFN15130_n_20599
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 247.09 0.0 247.118 0.163 ;
      END
   END FE_OFN15130_n_20599

   PIN FE_OFN15291_n_111917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.098 159.198 90.126 159.362 ;
      END
   END FE_OFN15291_n_111917

   PIN FE_OFN15295_n_111917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.562 159.198 128.59 159.362 ;
      END
   END FE_OFN15295_n_111917

   PIN FE_OFN15366_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 149.81 257.902 149.838 ;
      END
   END FE_OFN15366_delay_mul_ln34_unr5_unr5_stage2_stallmux_z_13_

   PIN FE_OFN15383_n_22225
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 240.498 0.0 240.526 0.163 ;
      END
   END FE_OFN15383_n_22225

   PIN FE_OFN15982_n_36821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.474 159.198 79.502 159.362 ;
      END
   END FE_OFN15982_n_36821

   PIN FE_OFN16234_n_40172
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 72.882 257.902 72.91 ;
      END
   END FE_OFN16234_n_40172

   PIN FE_OFN16237_n_40170
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 72.946 257.902 72.974 ;
      END
   END FE_OFN16237_n_40170

   PIN FE_OFN16239_n_40166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 72.882 257.902 72.91 ;
      END
   END FE_OFN16239_n_40166

   PIN FE_OFN16241_n_40166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 237.362 0.0 237.39 0.163 ;
      END
   END FE_OFN16241_n_40166

   PIN FE_OFN16256_n_40159
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 75.698 257.902 75.726 ;
      END
   END FE_OFN16256_n_40159

   PIN FE_OFN16649_n_7003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.53 0.0 228.558 0.163 ;
      END
   END FE_OFN16649_n_7003

   PIN FE_OFN17473_n_142961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 126.77 257.902 126.798 ;
      END
   END FE_OFN17473_n_142961

   PIN FE_OFN17490_n_142849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.866 159.198 106.894 159.362 ;
      END
   END FE_OFN17490_n_142849

   PIN FE_OFN17556_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.946 159.198 120.974 159.362 ;
      END
   END FE_OFN17556_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_

   PIN FE_OFN18570_b_4_7_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 138.29 0.163 138.318 ;
      END
   END FE_OFN18570_b_4_7_9

   PIN FE_OFN4555_n_142963
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.466 159.198 68.494 159.362 ;
      END
   END FE_OFN4555_n_142963

   PIN FE_OFN4568_n_41387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.538 159.198 151.566 159.362 ;
      END
   END FE_OFN4568_n_41387

   PIN FE_OFN4613_n_142796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.77 159.198 78.798 159.362 ;
      END
   END FE_OFN4613_n_142796

   PIN FE_OFN4646_n_142850
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.482 159.28 66.51 159.362 ;
      END
   END FE_OFN4646_n_142850

   PIN FE_OFN4665_n_137232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.962 159.198 86.99 159.362 ;
      END
   END FE_OFN4665_n_137232

   PIN FE_OFN4702_n_143619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.21 159.198 76.238 159.362 ;
      END
   END FE_OFN4702_n_143619

   PIN FE_OFN4762_n_137230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.242 159.198 80.27 159.362 ;
      END
   END FE_OFN4762_n_137230

   PIN FE_OFN4773_n_143004
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.61 159.198 82.638 159.362 ;
      END
   END FE_OFN4773_n_143004

   PIN FE_OFN4784_n_143003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.554 159.198 13.582 159.362 ;
      END
   END FE_OFN4784_n_143003

   PIN FE_OFN4791_n_41686
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 118.322 159.198 118.35 159.362 ;
      END
   END FE_OFN4791_n_41686

   PIN FE_OFN4796_n_143145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.122 159.198 75.15 159.362 ;
      END
   END FE_OFN4796_n_143145

   PIN FE_OFN4798_n_143146
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.002 159.198 94.03 159.362 ;
      END
   END FE_OFN4798_n_143146

   PIN FE_OFN4806_n_143143
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.698 159.198 123.726 159.362 ;
      END
   END FE_OFN4806_n_143143

   PIN FE_OFN4826_n_143199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.346 159.198 63.374 159.362 ;
      END
   END FE_OFN4826_n_143199

   PIN FE_OFN4885_n_36821
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.45 159.198 78.478 159.362 ;
      END
   END FE_OFN4885_n_36821

   PIN FE_OFN4999_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 157.362 257.902 157.39 ;
      END
   END FE_OFN4999_delay_mul_ln34_unr5_unr7_stage2_stallmux_z_11_

   PIN FE_OFN635_n_11194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 27.058 257.902 27.086 ;
      END
   END FE_OFN635_n_11194

   PIN FE_OFN637_n_8336
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.298 0.0 245.326 0.163 ;
      END
   END FE_OFN637_n_8336

   PIN FE_OFN654_n_8338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 244.082 0.0 244.11 0.163 ;
      END
   END FE_OFN654_n_8338

   PIN FE_OFN747_n_22238
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 167.09 0.0 167.118 0.163 ;
      END
   END FE_OFN747_n_22238

   PIN FE_OFN7582_n_40036
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.674 0.0 218.702 0.163 ;
      END
   END FE_OFN7582_n_40036

   PIN FE_OFN758_n_21703
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.346 0.0 199.374 0.163 ;
      END
   END FE_OFN758_n_21703

   PIN FE_OFN7819_n_40176
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 37.362 257.902 37.39 ;
      END
   END FE_OFN7819_n_40176

   PIN FE_OFN9214_delay_add_ln34_unr2_unr8_stage2_stallmux_q_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.186 0.0 67.214 0.163 ;
      END
   END FE_OFN9214_delay_add_ln34_unr2_unr8_stage2_stallmux_q_13_

   PIN FE_OFN9216_delay_add_ln34_unr2_unr8_stage2_stallmux_q_12_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.626 0.0 224.654 0.163 ;
      END
   END FE_OFN9216_delay_add_ln34_unr2_unr8_stage2_stallmux_q_12_

   PIN FE_OFN9895_b_4_7_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.674 159.198 74.702 159.362 ;
      END
   END FE_OFN9895_b_4_7_12

   PIN FE_OFN9897_b_4_7_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 72.434 159.198 72.462 159.362 ;
      END
   END FE_OFN9897_b_4_7_11

   PIN FE_OFN9899_b_4_7_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.354 159.198 90.382 159.362 ;
      END
   END FE_OFN9899_b_4_7_10

   PIN FE_OFN9905_b_4_7_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.578 159.198 70.606 159.362 ;
      END
   END FE_OFN9905_b_4_7_8

   PIN FE_OFN9908_b_4_7_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.994 159.198 75.022 159.362 ;
      END
   END FE_OFN9908_b_4_7_7

   PIN FE_OFN9910_b_4_7_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 75.058 159.198 75.086 159.362 ;
      END
   END FE_OFN9910_b_4_7_6

   PIN FE_OFN9911_b_4_7_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.994 159.198 75.022 159.362 ;
      END
   END FE_OFN9911_b_4_7_6

   PIN FE_OFN9913_b_4_7_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.674 159.198 82.702 159.362 ;
      END
   END FE_OFN9913_b_4_7_5

   PIN FE_OFN9914_b_4_7_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.13 159.198 86.158 159.362 ;
      END
   END FE_OFN9914_b_4_7_5

   PIN FE_OFN9916_b_4_7_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.514 159.198 78.542 159.362 ;
      END
   END FE_OFN9916_b_4_7_4

   PIN FE_OFN9917_b_4_7_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.41 159.198 95.438 159.362 ;
      END
   END FE_OFN9917_b_4_7_4

   PIN FE_OFN9919_b_4_7_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.738 159.198 82.766 159.362 ;
      END
   END FE_OFN9919_b_4_7_3

   PIN FE_OFN9920_b_4_7_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.706 159.198 86.734 159.362 ;
      END
   END FE_OFN9920_b_4_7_3

   PIN FE_OFN9922_b_4_7_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.602 159.198 87.63 159.362 ;
      END
   END FE_OFN9922_b_4_7_2

   PIN FE_OFN9923_b_4_7_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 101.81 159.198 101.838 159.362 ;
      END
   END FE_OFN9923_b_4_7_2

   PIN FE_OFN9925_b_4_7_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.994 159.198 51.022 159.362 ;
      END
   END FE_OFN9925_b_4_7_1

   PIN FE_OFN9928_b_4_7_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.786 159.198 76.814 159.362 ;
      END
   END FE_OFN9928_b_4_7_0

   PIN a_0_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.362 257.902 85.39 ;
      END
   END a_0_4_0

   PIN a_0_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.794 159.198 247.822 159.362 ;
      END
   END a_0_4_7

   PIN a_0_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 255.474 159.198 255.502 159.362 ;
      END
   END a_0_6_4

   PIN a_1_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.73 159.198 247.758 159.362 ;
      END
   END a_1_4_0

   PIN a_1_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.298 257.902 85.326 ;
      END
   END a_1_4_1

   PIN a_1_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.05 0.0 144.078 0.163 ;
      END
   END a_1_4_6

   PIN a_1_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 251.634 159.198 251.662 159.362 ;
      END
   END a_1_6_1

   PIN a_1_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 134.13 257.902 134.158 ;
      END
   END a_1_6_4

   PIN a_2_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 114.29 257.902 114.318 ;
      END
   END a_2_4_0

   PIN a_2_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 255.538 159.198 255.566 159.362 ;
      END
   END a_2_4_1

   PIN a_2_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 75.826 257.902 75.854 ;
      END
   END a_2_4_5

   PIN a_2_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 251.698 159.198 251.726 159.362 ;
      END
   END a_2_4_7

   PIN a_2_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.546 0.163 34.574 ;
      END
   END a_2_6_1

   PIN a_2_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 134.066 257.902 134.094 ;
      END
   END a_2_6_4

   PIN a_2_8_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 134.002 257.902 134.03 ;
      END
   END a_2_8_4

   PIN a_3_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 114.226 257.902 114.254 ;
      END
   END a_3_4_0

   PIN a_3_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 255.41 159.198 255.438 159.362 ;
      END
   END a_3_4_5

   PIN a_3_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.106 159.198 229.134 159.362 ;
      END
   END a_3_4_6

   PIN a_3_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 75.826 257.902 75.854 ;
      END
   END a_3_6_1

   PIN a_3_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 255.474 159.198 255.502 159.362 ;
      END
   END a_3_6_4

   PIN a_3_8_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 133.938 257.902 133.966 ;
      END
   END a_3_8_7

   PIN a_4_0_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 95.09 257.902 95.118 ;
      END
   END a_4_0_5

   PIN a_4_2_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.874 0.0 245.902 0.163 ;
      END
   END a_4_2_1

   PIN a_4_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 251.634 159.198 251.662 159.362 ;
      END
   END a_4_4_4

   PIN a_4_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 255.41 159.198 255.438 159.362 ;
      END
   END a_4_6_4

   PIN a_5_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.882 0.0 224.91 0.163 ;
      END
   END a_5_6_1

   PIN a_5_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 143.602 257.902 143.63 ;
      END
   END a_5_6_4

   PIN a_6_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 46.898 257.902 46.926 ;
      END
   END a_6_4_1

   PIN a_6_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 247.73 159.198 247.758 159.362 ;
      END
   END a_6_6_1

   PIN a_7_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 47.026 257.902 47.054 ;
      END
   END a_7_4_1

   PIN a_7_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 237.042 159.198 237.07 159.362 ;
      END
   END a_7_4_5

   PIN a_7_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 114.162 257.902 114.19 ;
      END
   END a_7_6_4

   PIN a_8_8_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 143.538 257.902 143.566 ;
      END
   END a_8_8_4

   PIN a_9_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 247.666 159.198 247.694 159.362 ;
      END
   END a_9_4_0

   PIN b_4_8_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 138.226 0.163 138.254 ;
      END
   END b_4_8_1

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.026 0.0 215.054 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_0_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.65 0.0 201.678 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_5_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 193.586 0.0 193.614 0.163 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_6_

   PIN delay_add_ln34_unr2_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 56.498 257.902 56.526 ;
      END
   END delay_add_ln34_unr2_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr3_unr0_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 91.954 257.902 91.982 ;
      END
   END delay_mul_ln34_unr3_unr0_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr3_unr5_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 153.778 257.902 153.806 ;
      END
   END delay_mul_ln34_unr3_unr5_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr3_unr7_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 99.762 257.902 99.79 ;
      END
   END delay_mul_ln34_unr3_unr7_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr3_unr7_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 198.962 0.0 198.99 0.163 ;
      END
   END delay_mul_ln34_unr3_unr7_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr3_unr7_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 80.498 257.902 80.526 ;
      END
   END delay_mul_ln34_unr3_unr7_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr3_unr8_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 88.114 257.902 88.142 ;
      END
   END delay_mul_ln34_unr3_unr8_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 201.65 159.198 201.678 159.362 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.29 159.198 90.318 159.362 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.226 159.198 90.254 159.362 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr4_unr0_stage2_stallmux_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.322 159.198 86.35 159.362 ;
      END
   END delay_mul_ln34_unr4_unr0_stage2_stallmux_z_7_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.29 159.198 242.318 159.362 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_q_15_

   PIN delay_mul_ln34_unr4_unr5_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.178 159.198 224.206 159.362 ;
      END
   END delay_mul_ln34_unr4_unr5_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.018 159.198 196.046 159.362 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_q_2_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 114.098 257.902 114.126 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 143.858 257.902 143.886 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 240.242 159.198 240.27 159.362 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr5_unr0_stage2_stallmux_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 124.338 257.902 124.366 ;
      END
   END delay_mul_ln34_unr5_unr0_stage2_stallmux_z_5_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 190.13 159.198 190.158 159.362 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_0_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 138.162 257.902 138.19 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_1_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 130.61 257.902 130.638 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_4_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_5_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 126.642 257.902 126.67 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_5_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 130.546 257.902 130.574 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr5_unr3_stage2_stallmux_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 107.506 257.902 107.534 ;
      END
   END delay_mul_ln34_unr5_unr3_stage2_stallmux_q_8_

   PIN delay_mul_ln34_unr5_unr5_stage2_stallmux_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.546 159.198 226.574 159.362 ;
      END
   END delay_mul_ln34_unr5_unr5_stage2_stallmux_z_10_

   PIN delay_mul_ln34_unr5_unr5_stage2_stallmux_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.162 159.198 186.19 159.362 ;
      END
   END delay_mul_ln34_unr5_unr5_stage2_stallmux_z_11_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 149.682 257.902 149.71 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_6_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 130.482 257.902 130.51 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_q_7_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 153.138 257.902 153.166 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_13_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 153.202 257.902 153.23 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_14_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 149.746 257.902 149.774 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_2_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 124.786 159.198 124.814 159.362 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_4_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_8_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 111.282 257.902 111.31 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_8_

   PIN delay_mul_ln34_unr5_unr7_stage2_stallmux_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 163.25 159.198 163.278 159.362 ;
      END
   END delay_mul_ln34_unr5_unr7_stage2_stallmux_z_9_

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 131.186 159.28 131.214 159.362 ;
      END
   END ispd_clk

   PIN mul_4646_72_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.386 159.198 78.414 159.362 ;
      END
   END mul_4646_72_n_116

   PIN mul_4646_72_n_124
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.154 159.198 63.182 159.362 ;
      END
   END mul_4646_72_n_124

   PIN mul_4646_72_n_212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.746 159.198 101.774 159.362 ;
      END
   END mul_4646_72_n_212

   PIN mul_4646_72_n_213
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.61 159.198 146.638 159.362 ;
      END
   END mul_4646_72_n_213

   PIN mul_4646_72_n_214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.922 159.198 143.95 159.362 ;
      END
   END mul_4646_72_n_214

   PIN mul_4646_72_n_96
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.386 159.198 86.414 159.362 ;
      END
   END mul_4646_72_n_96

   PIN mul_4646_72_n_97
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.49 0.0 101.518 0.163 ;
      END
   END mul_4646_72_n_97

   PIN mul_4646_72_n_98
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.554 0.0 101.582 0.163 ;
      END
   END mul_4646_72_n_98

   PIN mul_4650_72_n_288
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.546 159.198 58.574 159.362 ;
      END
   END mul_4650_72_n_288

   PIN mul_4650_72_n_307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.194 159.198 62.222 159.362 ;
      END
   END mul_4650_72_n_307

   PIN mul_4650_72_n_312
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.61 159.198 82.638 159.362 ;
      END
   END mul_4650_72_n_312

   PIN mul_4650_72_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.442 0.0 59.47 0.163 ;
      END
   END mul_4650_72_n_50

   PIN mul_4650_72_n_51
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.082 0.0 44.11 0.163 ;
      END
   END mul_4650_72_n_51

   PIN mul_4650_72_n_57
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.738 0.0 106.766 0.163 ;
      END
   END mul_4650_72_n_57

   PIN mul_4650_72_n_66
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.082 159.198 44.11 159.362 ;
      END
   END mul_4650_72_n_66

   PIN mul_4650_72_n_67
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.698 0.0 51.726 0.163 ;
      END
   END mul_4650_72_n_67

   PIN mul_4650_72_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.73 0.0 55.758 0.163 ;
      END
   END mul_4650_72_n_71

   PIN mul_4650_72_n_752
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.074 159.198 153.102 159.362 ;
      END
   END mul_4650_72_n_752

   PIN mul_4650_72_n_767
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.546 0.0 106.574 0.163 ;
      END
   END mul_4650_72_n_767

   PIN mul_4650_72_n_773
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.602 0.0 55.63 0.163 ;
      END
   END mul_4650_72_n_773

   PIN mul_4650_72_n_789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.914 0.0 36.942 0.163 ;
      END
   END mul_4650_72_n_789

   PIN mul_4650_72_n_837
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.426 0.0 61.454 0.163 ;
      END
   END mul_4650_72_n_837

   PIN mul_4650_72_n_840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.826 0.0 51.854 0.163 ;
      END
   END mul_4650_72_n_840

   PIN n_112253
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.53 159.198 36.558 159.362 ;
      END
   END n_112253

   PIN n_112259
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.418 159.198 146.446 159.362 ;
      END
   END n_112259

   PIN n_112755
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 136.434 159.198 136.462 159.362 ;
      END
   END n_112755

   PIN n_113329
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.218 159.198 103.246 159.362 ;
      END
   END n_113329

   PIN n_113795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.154 159.198 103.182 159.362 ;
      END
   END n_113795

   PIN n_113875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.61 0.0 82.638 0.163 ;
      END
   END n_113875

   PIN n_114487
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.418 159.198 82.446 159.362 ;
      END
   END n_114487

   PIN n_115523
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.89 159.198 51.918 159.362 ;
      END
   END n_115523

   PIN n_115564
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.266 159.198 113.294 159.362 ;
      END
   END n_115564

   PIN n_115565
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.618 159.198 117.646 159.362 ;
      END
   END n_115565

   PIN n_116610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.962 159.198 46.99 159.362 ;
      END
   END n_116610

   PIN n_116849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 113.266 159.198 113.294 159.362 ;
      END
   END n_116849

   PIN n_116850
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 113.202 159.198 113.23 159.362 ;
      END
   END n_116850

   PIN n_117661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.026 159.198 103.054 159.362 ;
      END
   END n_117661

   PIN n_117721
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.066 0.0 94.094 0.163 ;
      END
   END n_117721

   PIN n_119045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.786 159.198 28.814 159.362 ;
      END
   END n_119045

   PIN n_120348
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.986 159.198 48.014 159.362 ;
      END
   END n_120348

   PIN n_120860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.794 159.198 47.822 159.362 ;
      END
   END n_120860

   PIN n_121613
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.562 159.198 32.59 159.362 ;
      END
   END n_121613

   PIN n_121641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 124.85 159.198 124.878 159.362 ;
      END
   END n_121641

   PIN n_121888
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.554 0.0 69.582 0.163 ;
      END
   END n_121888

   PIN n_123339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.146 159.198 44.174 159.362 ;
      END
   END n_123339

   PIN n_124376
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.026 0.0 71.054 0.163 ;
      END
   END n_124376

   PIN n_124377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.49 0.0 69.518 0.163 ;
      END
   END n_124377

   PIN n_124389
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.546 159.198 74.574 159.362 ;
      END
   END n_124389

   PIN n_124393
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.746 0.0 93.774 0.163 ;
      END
   END n_124393

   PIN n_124629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.866 0.0 74.894 0.163 ;
      END
   END n_124629

   PIN n_124852
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.386 0.0 86.414 0.163 ;
      END
   END n_124852

   PIN n_124877
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.842 0.0 89.87 0.163 ;
      END
   END n_124877

   PIN n_125649
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.93 0.0 74.958 0.163 ;
      END
   END n_125649

   PIN n_126016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.306 159.198 32.334 159.362 ;
      END
   END n_126016

   PIN n_127097
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.834 0.0 78.862 0.163 ;
      END
   END n_127097

   PIN n_127103
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.866 0.0 66.894 0.163 ;
      END
   END n_127103

   PIN n_127612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.65 0.0 97.678 0.163 ;
      END
   END n_127612

   PIN n_128902
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.17 159.198 37.198 159.362 ;
      END
   END n_128902

   PIN n_129209
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 63.41 0.0 63.438 0.163 ;
      END
   END n_129209

   PIN n_129975
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 104.498 0.163 104.526 ;
      END
   END n_129975

   PIN n_133431
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.458 159.198 105.486 159.362 ;
      END
   END n_133431

   PIN n_134167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.274 0.0 44.302 0.163 ;
      END
   END n_134167

   PIN n_134694
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.762 0.0 51.79 0.163 ;
      END
   END n_134694

   PIN n_13477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.466 0.0 132.494 0.163 ;
      END
   END n_13477

   PIN n_13502
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 49.906 257.902 49.934 ;
      END
   END n_13502

   PIN n_137787
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 159.41 159.198 159.438 159.362 ;
      END
   END n_137787

   PIN n_137874
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 107.442 257.902 107.47 ;
      END
   END n_137874

   PIN n_143007
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.282 159.198 63.31 159.362 ;
      END
   END n_143007

   PIN n_144214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 42.226 257.902 42.254 ;
      END
   END n_144214

   PIN n_16610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.322 159.198 142.35 159.362 ;
      END
   END n_16610

   PIN n_16611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.514 159.198 142.542 159.362 ;
      END
   END n_16611

   PIN n_18394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.034 0.0 218.062 0.163 ;
      END
   END n_18394

   PIN n_18395
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 184.946 0.0 184.974 0.163 ;
      END
   END n_18395

   PIN n_18396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.586 0.0 201.614 0.163 ;
      END
   END n_18396

   PIN n_18397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.778 0.0 201.806 0.163 ;
      END
   END n_18397

   PIN n_18398
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 34.482 257.902 34.51 ;
      END
   END n_18398

   PIN n_18400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 34.546 257.902 34.574 ;
      END
   END n_18400

   PIN n_18779
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 189.746 0.0 189.774 0.163 ;
      END
   END n_18779

   PIN n_19896
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 7.986 257.902 8.014 ;
      END
   END n_19896

   PIN n_19897
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 234.802 0.0 234.83 0.163 ;
      END
   END n_19897

   PIN n_19898
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 174.834 0.0 174.862 0.163 ;
      END
   END n_19898

   PIN n_19899
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.514 0.0 182.542 0.163 ;
      END
   END n_19899

   PIN n_20359
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.466 0.0 228.494 0.163 ;
      END
   END n_20359

   PIN n_20449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 151.73 159.198 151.758 159.362 ;
      END
   END n_20449

   PIN n_20564
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.93 0.0 170.958 0.163 ;
      END
   END n_20564

   PIN n_20565
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.186 0.0 163.214 0.163 ;
      END
   END n_20565

   PIN n_20644
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 30.706 257.902 30.734 ;
      END
   END n_20644

   PIN n_20800
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 236.21 0.0 236.238 0.163 ;
      END
   END n_20800

   PIN n_21064
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.018 159.198 148.046 159.362 ;
      END
   END n_21064

   PIN n_21065
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.05 159.198 176.078 159.362 ;
      END
   END n_21065

   PIN n_21066
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.826 159.198 211.854 159.362 ;
      END
   END n_21066

   PIN n_21069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 167.09 159.198 167.118 159.362 ;
      END
   END n_21069

   PIN n_21096
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 66.29 257.902 66.318 ;
      END
   END n_21096

   PIN n_21097
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 66.226 257.902 66.254 ;
      END
   END n_21097

   PIN n_21145
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.802 0.0 170.83 0.163 ;
      END
   END n_21145

   PIN n_21358
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 142.386 159.198 142.414 159.362 ;
      END
   END n_21358

   PIN n_21365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 66.354 257.902 66.382 ;
      END
   END n_21365

   PIN n_21400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.954 159.198 147.982 159.362 ;
      END
   END n_21400

   PIN n_21449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.466 159.198 164.494 159.362 ;
      END
   END n_21449

   PIN n_21451
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 236.146 0.0 236.174 0.163 ;
      END
   END n_21451

   PIN n_21616
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.81 0.0 197.838 0.163 ;
      END
   END n_21616

   PIN n_21617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.746 0.0 197.774 0.163 ;
      END
   END n_21617

   PIN n_21621
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.458 0.0 201.486 0.163 ;
      END
   END n_21621

   PIN n_21671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 240.05 0.0 240.078 0.163 ;
      END
   END n_21671

   PIN n_21890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 197.682 0.0 197.71 0.163 ;
      END
   END n_21890

   PIN n_22137
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.746 159.198 205.774 159.362 ;
      END
   END n_22137

   PIN n_22166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.362 0.0 205.39 0.163 ;
      END
   END n_22166

   PIN n_22167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 209.33 0.0 209.358 0.163 ;
      END
   END n_22167

   PIN n_22235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.866 0.0 170.894 0.163 ;
      END
   END n_22235

   PIN n_22448
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 72.754 257.902 72.782 ;
      END
   END n_22448

   PIN n_22449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 61.426 257.902 61.454 ;
      END
   END n_22449

   PIN n_22475
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.714 0.0 201.742 0.163 ;
      END
   END n_22475

   PIN n_22476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 201.65 0.0 201.678 0.163 ;
      END
   END n_22476

   PIN n_22516
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.49 0.0 205.518 0.163 ;
      END
   END n_22516

   PIN n_22541
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.426 0.0 205.454 0.163 ;
      END
   END n_22541

   PIN n_22817
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.21 0.0 172.238 0.163 ;
      END
   END n_22817

   PIN n_23018
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 37.298 257.902 37.326 ;
      END
   END n_23018

   PIN n_23041
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.146 0.0 140.174 0.163 ;
      END
   END n_23041

   PIN n_23125
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 104.498 257.902 104.526 ;
      END
   END n_23125

   PIN n_23330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 99.826 257.902 99.854 ;
      END
   END n_23330

   PIN n_23555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 132.53 0.0 132.558 0.163 ;
      END
   END n_23555

   PIN n_23647
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 94.962 257.902 94.99 ;
      END
   END n_23647

   PIN n_23667
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.026 0.0 119.054 0.163 ;
      END
   END n_23667

   PIN n_23669
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 105.458 0.0 105.486 0.163 ;
      END
   END n_23669

   PIN n_23722
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 105.586 0.0 105.614 0.163 ;
      END
   END n_23722

   PIN n_23768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 118.962 257.902 118.99 ;
      END
   END n_23768

   PIN n_24318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.234 0.0 117.262 0.163 ;
      END
   END n_24318

   PIN n_24395
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.714 159.198 201.742 159.362 ;
      END
   END n_24395

   PIN n_24709
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.522 0.0 201.55 0.163 ;
      END
   END n_24709

   PIN n_25046
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 94.898 257.902 94.926 ;
      END
   END n_25046

   PIN n_26039
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.026 0.0 207.054 0.163 ;
      END
   END n_26039

   PIN n_26266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 104.626 257.902 104.654 ;
      END
   END n_26266

   PIN n_26268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 57.522 257.902 57.55 ;
      END
   END n_26268

   PIN n_26406
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.674 159.198 218.702 159.362 ;
      END
   END n_26406

   PIN n_26895
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 85.746 257.902 85.774 ;
      END
   END n_26895

   PIN n_26897
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 69.106 257.902 69.134 ;
      END
   END n_26897

   PIN n_26908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 27.314 257.902 27.342 ;
      END
   END n_26908

   PIN n_27622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.946 159.198 216.974 159.362 ;
      END
   END n_27622

   PIN n_27970
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.45 0.0 182.478 0.163 ;
      END
   END n_27970

   PIN n_27972
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.386 0.0 182.414 0.163 ;
      END
   END n_27972

   PIN n_2799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.466 0.0 36.494 0.163 ;
      END
   END n_2799

   PIN n_28572
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.554 159.198 205.582 159.362 ;
      END
   END n_28572

   PIN n_28574
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.386 159.198 230.414 159.362 ;
      END
   END n_28574

   PIN n_2861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 170.93 159.198 170.958 159.362 ;
      END
   END n_2861

   PIN n_2871
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.674 0.0 138.702 0.163 ;
      END
   END n_2871

   PIN n_28733
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.258 159.198 230.286 159.362 ;
      END
   END n_28733

   PIN n_29056
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.634 159.198 227.662 159.362 ;
      END
   END n_29056

   PIN n_29058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 227.442 159.198 227.47 159.362 ;
      END
   END n_29058

   PIN n_32114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.37 159.198 80.398 159.362 ;
      END
   END n_32114

   PIN n_32115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 80.178 159.198 80.206 159.362 ;
      END
   END n_32115

   PIN n_32440
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.898 159.198 86.926 159.362 ;
      END
   END n_32440

   PIN n_32718
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.322 159.198 38.35 159.362 ;
      END
   END n_32718

   PIN n_32740
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.442 159.198 51.47 159.362 ;
      END
   END n_32740

   PIN n_32741
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.25 159.198 51.278 159.362 ;
      END
   END n_32741

   PIN n_32769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.682 159.198 69.71 159.362 ;
      END
   END n_32769

   PIN n_33082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.746 159.198 61.774 159.362 ;
      END
   END n_33082

   PIN n_33167
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.018 159.198 44.046 159.362 ;
      END
   END n_33167

   PIN n_33364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.354 159.198 82.382 159.362 ;
      END
   END n_33364

   PIN n_33881
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.258 159.198 86.286 159.362 ;
      END
   END n_33881

   PIN n_34014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.306 159.198 40.334 159.362 ;
      END
   END n_34014

   PIN n_34377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 40.242 159.198 40.27 159.362 ;
      END
   END n_34377

   PIN n_34609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.306 159.198 80.334 159.362 ;
      END
   END n_34609

   PIN n_34610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.498 159.198 80.526 159.362 ;
      END
   END n_34610

   PIN n_34731
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.194 159.198 86.222 159.362 ;
      END
   END n_34731

   PIN n_34808
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.506 159.198 3.534 159.362 ;
      END
   END n_34808

   PIN n_3513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 171.058 159.198 171.086 159.362 ;
      END
   END n_3513

   PIN n_35434
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.834 159.198 54.862 159.362 ;
      END
   END n_35434

   PIN n_36613
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.218 159.198 63.246 159.362 ;
      END
   END n_36613

   PIN n_37477
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.394 159.198 25.422 159.362 ;
      END
   END n_37477

   PIN n_37556
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.554 159.198 101.582 159.362 ;
      END
   END n_37556

   PIN n_37622
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.634 159.198 91.662 159.362 ;
      END
   END n_37622

   PIN n_37665
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.202 159.198 145.23 159.362 ;
      END
   END n_37665

   PIN n_37690
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.802 159.198 74.83 159.362 ;
      END
   END n_37690

   PIN n_382
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 152.882 159.198 152.91 159.362 ;
      END
   END n_382

   PIN n_39240
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.042 159.198 69.07 159.362 ;
      END
   END n_39240

   PIN n_39453
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.81 0.0 101.838 0.163 ;
      END
   END n_39453

   PIN n_39845
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.306 159.198 136.334 159.362 ;
      END
   END n_39845

   PIN n_40155
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.821 27.186 257.902 27.214 ;
      END
   END n_40155

   PIN n_40158
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 80.69 257.902 80.718 ;
      END
   END n_40158

   PIN n_40330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 72.818 257.902 72.846 ;
      END
   END n_40330

   PIN n_40445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 56.562 257.902 56.59 ;
      END
   END n_40445

   PIN n_40476
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 73.074 257.902 73.102 ;
      END
   END n_40476

   PIN n_40561
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 92.146 257.902 92.174 ;
      END
   END n_40561

   PIN n_40564
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 88.242 257.902 88.27 ;
      END
   END n_40564

   PIN n_40626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 75.762 257.902 75.79 ;
      END
   END n_40626

   PIN n_40648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 75.698 257.902 75.726 ;
      END
   END n_40648

   PIN n_40695
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 202.738 0.0 202.766 0.163 ;
      END
   END n_40695

   PIN n_40706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 75.762 257.902 75.79 ;
      END
   END n_40706

   PIN n_40727
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 88.306 257.902 88.334 ;
      END
   END n_40727

   PIN n_48178
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.098 159.198 74.126 159.362 ;
      END
   END n_48178

   PIN n_48510
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.122 159.198 67.15 159.362 ;
      END
   END n_48510

   PIN n_48907
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.49 159.198 77.518 159.362 ;
      END
   END n_48907

   PIN n_49236
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 66.162 257.902 66.19 ;
      END
   END n_49236

   PIN n_5058
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.642 0.0 150.67 0.163 ;
      END
   END n_5058

   PIN n_5059
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 150.834 0.0 150.862 0.163 ;
      END
   END n_5059

   PIN n_5115
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 147.762 159.198 147.79 159.362 ;
      END
   END n_5115

   PIN n_51768
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.738 159.198 74.766 159.362 ;
      END
   END n_51768

   PIN n_54235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.426 159.198 77.454 159.362 ;
      END
   END n_54235

   PIN n_54706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 66.098 257.902 66.126 ;
      END
   END n_54706

   PIN n_5505
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.37 159.198 136.398 159.362 ;
      END
   END n_5505

   PIN n_5571
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 162.994 0.0 163.022 0.163 ;
      END
   END n_5571

   PIN n_57100
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.298 159.198 77.326 159.362 ;
      END
   END n_57100

   PIN n_58492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 72.818 257.902 72.846 ;
      END
   END n_58492

   PIN n_58941
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.498 159.198 72.526 159.362 ;
      END
   END n_58941

   PIN n_60391
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 76.658 257.902 76.686 ;
      END
   END n_60391

   PIN n_6364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.994 159.198 171.022 159.362 ;
      END
   END n_6364

   PIN n_63870
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 257.739 80.498 257.902 80.526 ;
      END
   END n_63870

   PIN n_6635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 257.739 153.138 257.902 153.166 ;
      END
   END n_6635

   PIN n_7003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.962 0.0 246.99 0.163 ;
      END
   END n_7003

   PIN n_7337
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.194 159.198 94.222 159.362 ;
      END
   END n_7337

   PIN n_7696
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.114 0.0 48.142 0.163 ;
      END
   END n_7696

   PIN n_7848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 94.13 159.198 94.158 159.362 ;
      END
   END n_7848

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 257.902 159.362 ;
      LAYER V1 ;
         RECT 0.0 0.0 257.902 159.362 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 257.902 159.362 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 257.902 159.362 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 257.902 159.362 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 257.902 159.362 ;
      LAYER M1 ;
         RECT 0.0 0.0 257.902 159.362 ;
   END
END h1_mgc_matrix_mult_b

MACRO h0_mgc_matrix_mult_b
   CLASS BLOCK ;
   FOREIGN h0 ;
   ORIGIN 0 0 ;
   SIZE 313.394 BY 122.24 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN10233_b_2_6_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 86.258 0.163 86.286 ;
      END
   END FE_OFN10233_b_2_6_0

   PIN FE_OFN10257_b_2_4_6
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.714 0.163 97.742 ;
      END
   END FE_OFN10257_b_2_4_6

   PIN FE_OFN10260_b_2_4_5
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.37 122.077 136.398 122.24 ;
      END
   END FE_OFN10260_b_2_4_5

   PIN FE_OFN10293_b_2_2_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.33 0.163 113.358 ;
      END
   END FE_OFN10293_b_2_2_3

   PIN FE_OFN1071_n_16034
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 284.018 122.077 284.046 122.24 ;
      END
   END FE_OFN1071_n_16034

   PIN FE_OFN1086_n_21187
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.386 122.077 238.414 122.24 ;
      END
   END FE_OFN1086_n_21187

   PIN FE_OFN11430_n_142905
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 90.226 0.163 90.254 ;
      END
   END FE_OFN11430_n_142905

   PIN FE_OFN11434_n_142919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.81 0.163 101.838 ;
      END
   END FE_OFN11434_n_142919

   PIN FE_OFN11435_n_142919
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 211.378 122.077 211.406 122.24 ;
      END
   END FE_OFN11435_n_142919

   PIN FE_OFN1157_n_10648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.602 122.077 215.63 122.24 ;
      END
   END FE_OFN1157_n_10648

   PIN FE_OFN11706_n_142947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.45 0.163 118.478 ;
      END
   END FE_OFN11706_n_142947

   PIN FE_OFN11707_n_142947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.802 0.163 82.83 ;
      END
   END FE_OFN11707_n_142947

   PIN FE_OFN12301_n_111727
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.458 122.077 153.486 122.24 ;
      END
   END FE_OFN12301_n_111727

   PIN FE_OFN12386_n_142906
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.874 122.077 45.902 122.24 ;
      END
   END FE_OFN12386_n_142906

   PIN FE_OFN12400_n_694
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.842 0.163 113.87 ;
      END
   END FE_OFN12400_n_694

   PIN FE_OFN12617_n_112689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.778 122.077 137.806 122.24 ;
      END
   END FE_OFN12617_n_112689

   PIN FE_OFN12618_n_112689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 133.746 122.077 133.774 122.24 ;
      END
   END FE_OFN12618_n_112689

   PIN FE_OFN13018_n_142950
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 97.842 0.163 97.87 ;
      END
   END FE_OFN13018_n_142950

   PIN FE_OFN15062_n_12711
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.29 122.077 34.318 122.24 ;
      END
   END FE_OFN15062_n_12711

   PIN FE_OFN15077_n_14458
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 214.642 122.077 214.67 122.24 ;
      END
   END FE_OFN15077_n_14458

   PIN FE_OFN15252_n_39084
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.514 0.163 118.542 ;
      END
   END FE_OFN15252_n_39084

   PIN FE_OFN15923_n_143045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.93 0.163 74.958 ;
      END
   END FE_OFN15923_n_143045

   PIN FE_OFN15925_n_112550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.978 122.077 5.006 122.24 ;
      END
   END FE_OFN15925_n_112550

   PIN FE_OFN15930_n_143241
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.482 0.163 98.51 ;
      END
   END FE_OFN15930_n_143241

   PIN FE_OFN16294_delay_add_ln34_unr2_unr3_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.066 122.077 134.094 122.24 ;
      END
   END FE_OFN16294_delay_add_ln34_unr2_unr3_stage2_stallmux_q_15_

   PIN FE_OFN16366_b_2_4_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.218 122.077 119.246 122.24 ;
      END
   END FE_OFN16366_b_2_4_1

   PIN FE_OFN16771_n_16098
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 237.938 122.077 237.966 122.24 ;
      END
   END FE_OFN16771_n_16098

   PIN FE_OFN17162_n_132699
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.778 0.163 105.806 ;
      END
   END FE_OFN17162_n_132699

   PIN FE_OFN17165_n_134675
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.466 122.077 172.494 122.24 ;
      END
   END FE_OFN17165_n_134675

   PIN FE_OFN17200_n_16166
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 206.962 122.077 206.99 122.24 ;
      END
   END FE_OFN17200_n_16166

   PIN FE_OFN17265_n_140245
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 105.778 0.163 105.806 ;
      END
   END FE_OFN17265_n_140245

   PIN FE_OFN18609_b_2_2_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.522 0.163 113.55 ;
      END
   END FE_OFN18609_b_2_2_0

   PIN FE_OFN18810_n_143645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.298 0.163 109.326 ;
      END
   END FE_OFN18810_n_143645

   PIN FE_OFN19059_n_19681
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 110.258 0.163 110.286 ;
      END
   END FE_OFN19059_n_19681

   PIN FE_OFN19145_n_143045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.642 0.163 78.67 ;
      END
   END FE_OFN19145_n_143045

   PIN FE_OFN19307_b_2_2_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.714 122.077 49.742 122.24 ;
      END
   END FE_OFN19307_b_2_2_1

   PIN FE_OFN2160_n_19626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 214.77 122.077 214.798 122.24 ;
      END
   END FE_OFN2160_n_19626

   PIN FE_OFN2283_n_19629
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.826 122.077 91.854 122.24 ;
      END
   END FE_OFN2283_n_19629

   PIN FE_OFN3286_n_117368
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.05 122.077 88.078 122.24 ;
      END
   END FE_OFN3286_n_117368

   PIN FE_OFN3294_n_8246
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 239.41 122.077 239.438 122.24 ;
      END
   END FE_OFN3294_n_8246

   PIN FE_OFN3442_n_12341
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 216.562 122.077 216.59 122.24 ;
      END
   END FE_OFN3442_n_12341

   PIN FE_OFN3574_n_133235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.906 0.163 97.934 ;
      END
   END FE_OFN3574_n_133235

   PIN FE_OFN3613_n_112427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.122 122.077 123.15 122.24 ;
      END
   END FE_OFN3613_n_112427

   PIN FE_OFN3656_n_112550
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 85.49 0.163 85.518 ;
      END
   END FE_OFN3656_n_112550

   PIN FE_OFN3723_n_143241
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.658 122.077 100.686 122.24 ;
      END
   END FE_OFN3723_n_143241

   PIN FE_OFN606_n_8387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.842 122.077 145.87 122.24 ;
      END
   END FE_OFN606_n_8387

   PIN FE_OFN703_n_21657
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 236.466 122.077 236.494 122.24 ;
      END
   END FE_OFN703_n_21657

   PIN FE_OFN757_n_21703
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 214.002 122.077 214.03 122.24 ;
      END
   END FE_OFN757_n_21703

   PIN FE_OFN797_n_21129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 237.874 122.077 237.902 122.24 ;
      END
   END FE_OFN797_n_21129

   PIN add_5900_51_n_148
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 264.818 122.077 264.846 122.24 ;
      END
   END add_5900_51_n_148

   PIN add_5900_51_n_77
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.146 122.077 180.174 122.24 ;
      END
   END add_5900_51_n_77

   PIN delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.77 122.077 118.798 122.24 ;
      END
   END delay_add_ln34_unr2_unr1_stage2_stallmux_q_15_

   PIN delay_add_ln34_unr2_unr2_stage2_stallmux_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 149.554 122.077 149.582 122.24 ;
      END
   END delay_add_ln34_unr2_unr2_stage2_stallmux_z_12_

   PIN delay_add_ln34_unr2_unr3_stage2_stallmux_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 203.378 122.077 203.406 122.24 ;
      END
   END delay_add_ln34_unr2_unr3_stage2_stallmux_q_10_

   PIN delay_add_ln34_unr2_unr3_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 141.81 122.077 141.838 122.24 ;
      END
   END delay_add_ln34_unr2_unr3_stage2_stallmux_q_3_

   PIN delay_add_ln34_unr2_unr3_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 224.882 122.077 224.91 122.24 ;
      END
   END delay_add_ln34_unr2_unr3_stage2_stallmux_q_4_

   PIN delay_add_ln34_unr2_unr3_stage2_stallmux_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.29 122.077 130.318 122.24 ;
      END
   END delay_add_ln34_unr2_unr3_stage2_stallmux_q_8_

   PIN delay_add_ln34_unr2_unr5_stage2_stallmux_q_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.482 122.077 122.51 122.24 ;
      END
   END delay_add_ln34_unr2_unr5_stage2_stallmux_q_14_

   PIN delay_add_ln34_unr2_unr5_stage2_stallmux_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.586 122.077 145.614 122.24 ;
      END
   END delay_add_ln34_unr2_unr5_stage2_stallmux_q_7_

   PIN delay_add_ln34_unr2_unr5_stage2_stallmux_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.106 122.077 205.134 122.24 ;
      END
   END delay_add_ln34_unr2_unr5_stage2_stallmux_q_8_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 134.066 122.077 134.094 122.24 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_3_

   PIN delay_add_ln34_unr2_unr7_stage2_stallmux_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.282 122.077 191.31 122.24 ;
      END
   END delay_add_ln34_unr2_unr7_stage2_stallmux_q_4_

   PIN delay_add_ln34_unr2_unr8_stage2_stallmux_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 210.93 122.077 210.958 122.24 ;
      END
   END delay_add_ln34_unr2_unr8_stage2_stallmux_q_3_

   PIN mul_4665_72_n_202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.362 0.163 117.39 ;
      END
   END mul_4665_72_n_202

   PIN mul_4665_72_n_221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.146 122.077 28.174 122.24 ;
      END
   END mul_4665_72_n_221

   PIN mul_4665_72_n_230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.578 122.077 30.606 122.24 ;
      END
   END mul_4665_72_n_230

   PIN mul_4665_72_n_295
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.362 0.163 109.39 ;
      END
   END mul_4665_72_n_295

   PIN mul_4665_72_n_337
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 89.97 0.163 89.998 ;
      END
   END mul_4665_72_n_337

   PIN mul_4665_72_n_848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.074 0.163 105.102 ;
      END
   END mul_4665_72_n_848

   PIN mul_4667_72_n_184
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.218 122.077 111.246 122.24 ;
      END
   END mul_4667_72_n_184

   PIN mul_4667_72_n_265
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 26.61 122.077 26.638 122.24 ;
      END
   END mul_4667_72_n_265

   PIN mul_4667_72_n_304
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.162 0.163 98.19 ;
      END
   END mul_4667_72_n_304

   PIN mul_4667_72_n_308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.45 0.163 86.478 ;
      END
   END mul_4667_72_n_308

   PIN mul_4667_72_n_316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.138 122.077 65.166 122.24 ;
      END
   END mul_4667_72_n_316

   PIN mul_4667_72_n_323
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.858 122.077 79.886 122.24 ;
      END
   END mul_4667_72_n_323

   PIN mul_4667_72_n_324
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.738 122.077 82.766 122.24 ;
      END
   END mul_4667_72_n_324

   PIN mul_4667_72_n_327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.874 0.163 101.902 ;
      END
   END mul_4667_72_n_327

   PIN mul_4667_72_n_66
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.698 122.077 3.726 122.24 ;
      END
   END mul_4667_72_n_66

   PIN mul_4669_72_n_225
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.37 0.163 40.398 ;
      END
   END mul_4669_72_n_225

   PIN mul_4669_72_n_304
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.706 0.163 78.734 ;
      END
   END mul_4669_72_n_304

   PIN mul_4669_72_n_314
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.258 0.163 102.286 ;
      END
   END mul_4669_72_n_314

   PIN mul_4669_72_n_316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.194 0.163 102.222 ;
      END
   END mul_4669_72_n_316

   PIN mul_4669_72_n_66
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.186 0.163 67.214 ;
      END
   END mul_4669_72_n_66

   PIN mul_ln34_unr0_unr6_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.354 122.077 130.382 122.24 ;
      END
   END mul_ln34_unr0_unr6_z_14_

   PIN mul_ln34_unr2_unr2_z_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.426 122.077 149.454 122.24 ;
      END
   END mul_ln34_unr2_unr2_z_0_

   PIN mul_ln34_unr2_unr2_z_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 264.818 122.077 264.846 122.24 ;
      END
   END mul_ln34_unr2_unr2_z_14_

   PIN mul_ln34_unr2_unr2_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.786 122.077 164.814 122.24 ;
      END
   END mul_ln34_unr2_unr2_z_7_

   PIN n_10378
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.794 122.077 95.822 122.24 ;
      END
   END n_10378

   PIN n_10669
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.306 122.077 128.334 122.24 ;
      END
   END n_10669

   PIN n_11011
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.666 122.077 7.694 122.24 ;
      END
   END n_11011

   PIN n_111968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.09 122.077 15.118 122.24 ;
      END
   END n_111968

   PIN n_112778
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 113.266 313.394 113.294 ;
      END
   END n_112778

   PIN n_112779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 55.858 313.394 55.886 ;
      END
   END n_112779

   PIN n_112812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 67.25 313.394 67.278 ;
      END
   END n_112812

   PIN n_112817
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 101.554 0.163 101.582 ;
      END
   END n_112817

   PIN n_112831
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 312.37 122.077 312.398 122.24 ;
      END
   END n_112831

   PIN n_112845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 295.666 122.077 295.694 122.24 ;
      END
   END n_112845

   PIN n_112880
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 254.514 122.077 254.542 122.24 ;
      END
   END n_112880

   PIN n_112890
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.546 0.163 82.574 ;
      END
   END n_112890

   PIN n_112959
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.682 0.163 109.71 ;
      END
   END n_112959

   PIN n_113054
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 241.714 122.077 241.742 122.24 ;
      END
   END n_113054

   PIN n_113100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.042 0.163 109.07 ;
      END
   END n_113100

   PIN n_113160
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 110.13 0.163 110.158 ;
      END
   END n_113160

   PIN n_113191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 106.098 0.163 106.126 ;
      END
   END n_113191

   PIN n_113195
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 44.978 313.394 45.006 ;
      END
   END n_113195

   PIN n_113217
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.57 122.077 307.598 122.24 ;
      END
   END n_113217

   PIN n_113223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.866 0.163 82.894 ;
      END
   END n_113223

   PIN n_113308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 85.554 0.163 85.582 ;
      END
   END n_113308

   PIN n_113317
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 85.298 0.163 85.326 ;
      END
   END n_113317

   PIN n_113342
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.61 122.077 26.638 122.24 ;
      END
   END n_113342

   PIN n_113343
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.674 122.077 26.702 122.24 ;
      END
   END n_113343

   PIN n_113447
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 163.506 122.077 163.534 122.24 ;
      END
   END n_113447

   PIN n_113479
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.522 122.077 241.55 122.24 ;
      END
   END n_113479

   PIN n_113480
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.138 0.163 105.166 ;
      END
   END n_113480

   PIN n_113481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.202 0.163 105.23 ;
      END
   END n_113481

   PIN n_113503
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.106 122.077 5.134 122.24 ;
      END
   END n_113503

   PIN n_113516
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.738 122.077 26.766 122.24 ;
      END
   END n_113516

   PIN n_113517
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.802 122.077 26.83 122.24 ;
      END
   END n_113517

   PIN n_113545
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 106.162 0.163 106.19 ;
      END
   END n_113545

   PIN n_113830
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 299.25 122.077 299.278 122.24 ;
      END
   END n_113830

   PIN n_113933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.01 122.077 161.038 122.24 ;
      END
   END n_113933

   PIN n_113934
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.882 122.077 160.91 122.24 ;
      END
   END n_113934

   PIN n_114134
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 74.93 0.163 74.958 ;
      END
   END n_114134

   PIN n_114136
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.586 0.163 113.614 ;
      END
   END n_114136

   PIN n_114331
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 78.834 0.163 78.862 ;
      END
   END n_114331

   PIN n_114597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.946 122.077 160.974 122.24 ;
      END
   END n_114597

   PIN n_114598
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 161.202 122.077 161.23 122.24 ;
      END
   END n_114598

   PIN n_114821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.97 0.163 97.998 ;
      END
   END n_114821

   PIN n_114951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 63.41 0.163 63.438 ;
      END
   END n_114951

   PIN n_115117
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 110.322 0.163 110.35 ;
      END
   END n_115117

   PIN n_115119
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.122 0.163 75.15 ;
      END
   END n_115119

   PIN n_115219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.514 0.163 86.542 ;
      END
   END n_115219

   PIN n_116269
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.298 0.163 69.326 ;
      END
   END n_116269

   PIN n_116470
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.602 122.077 7.63 122.24 ;
      END
   END n_116470

   PIN n_117525
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.986 122.077 312.014 122.24 ;
      END
   END n_117525

   PIN n_117559
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 303.154 122.077 303.182 122.24 ;
      END
   END n_117559

   PIN n_117560
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 312.05 122.077 312.078 122.24 ;
      END
   END n_117560

   PIN n_117582
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 93.682 0.163 93.71 ;
      END
   END n_117582

   PIN n_117603
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.906 0.163 113.934 ;
      END
   END n_117603

   PIN n_117620
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.61 0.163 82.638 ;
      END
   END n_117620

   PIN n_118017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.106 0.163 109.134 ;
      END
   END n_118017

   PIN n_118035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 299.378 122.077 299.406 122.24 ;
      END
   END n_118035

   PIN n_118166
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.146 122.077 84.174 122.24 ;
      END
   END n_118166

   PIN n_118364
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 5.042 122.077 5.07 122.24 ;
      END
   END n_118364

   PIN n_119552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.266 0.163 105.294 ;
      END
   END n_119552

   PIN n_119619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 222.322 122.077 222.35 122.24 ;
      END
   END n_119619

   PIN n_119690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.034 0.163 114.062 ;
      END
   END n_119690

   PIN n_119691
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 117.618 0.163 117.646 ;
      END
   END n_119691

   PIN n_119709
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.226 0.163 114.254 ;
      END
   END n_119709

   PIN n_119812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.834 122.077 22.862 122.24 ;
      END
   END n_119812

   PIN n_119886
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 233.01 122.077 233.038 122.24 ;
      END
   END n_119886

   PIN n_119969
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 97.906 0.163 97.934 ;
      END
   END n_119969

   PIN n_120042
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.842 0.163 105.87 ;
      END
   END n_120042

   PIN n_120044
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 85.362 0.163 85.39 ;
      END
   END n_120044

   PIN n_120045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.65 0.163 113.678 ;
      END
   END n_120045

   PIN n_120129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.994 0.163 75.022 ;
      END
   END n_120129

   PIN n_120131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.362 0.163 69.39 ;
      END
   END n_120131

   PIN n_120499
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.29 0.163 90.318 ;
      END
   END n_120499

   PIN n_120794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.778 0.163 97.806 ;
      END
   END n_120794

   PIN n_121083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.81 0.163 117.838 ;
      END
   END n_121083

   PIN n_121084
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.81 0.163 109.838 ;
      END
   END n_121084

   PIN n_121196
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 312.434 122.077 312.462 122.24 ;
      END
   END n_121196

   PIN n_121291
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 307.058 122.077 307.086 122.24 ;
      END
   END n_121291

   PIN n_121522
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 253.17 122.077 253.198 122.24 ;
      END
   END n_121522

   PIN n_121732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 287.794 122.077 287.822 122.24 ;
      END
   END n_121732

   PIN n_121779
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.978 0.163 61.006 ;
      END
   END n_121779

   PIN n_121908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.746 0.163 93.774 ;
      END
   END n_121908

   PIN n_121917
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.418 0.163 82.446 ;
      END
   END n_121917

   PIN n_121918
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.674 0.163 82.702 ;
      END
   END n_121918

   PIN n_122005
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.122 122.077 107.15 122.24 ;
      END
   END n_122005

   PIN n_122026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 94.002 0.163 94.03 ;
      END
   END n_122026

   PIN n_122106
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.386 0.163 94.414 ;
      END
   END n_122106

   PIN n_122300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.21 122.077 84.238 122.24 ;
      END
   END n_122300

   PIN n_122476
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.33 122.077 153.358 122.24 ;
      END
   END n_122476

   PIN n_122532
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 237.81 122.077 237.838 122.24 ;
      END
   END n_122532

   PIN n_123300
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 69.426 0.163 69.454 ;
      END
   END n_123300

   PIN n_123316
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 97.778 0.163 97.806 ;
      END
   END n_123316

   PIN n_123618
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.466 122.077 84.494 122.24 ;
      END
   END n_123618

   PIN n_123955
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 312.498 122.077 312.526 122.24 ;
      END
   END n_123955

   PIN n_124058
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.73 0.163 55.758 ;
      END
   END n_124058

   PIN n_124589
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 11.314 122.077 11.342 122.24 ;
      END
   END n_124589

   PIN n_124590
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.378 122.077 11.406 122.24 ;
      END
   END n_124590

   PIN n_124859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 247.602 122.077 247.63 122.24 ;
      END
   END n_124859

   PIN n_125049
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 101.81 313.394 101.838 ;
      END
   END n_125049

   PIN n_125190
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 257.074 122.077 257.102 122.24 ;
      END
   END n_125190

   PIN n_125260
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 86.578 313.394 86.606 ;
      END
   END n_125260

   PIN n_125261
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.634 122.077 307.662 122.24 ;
      END
   END n_125261

   PIN n_125371
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.322 0.163 94.35 ;
      END
   END n_125371

   PIN n_125378
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.642 0.163 94.67 ;
      END
   END n_125378

   PIN n_125536
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.506 122.077 235.534 122.24 ;
      END
   END n_125536

   PIN n_125537
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 231.538 122.077 231.566 122.24 ;
      END
   END n_125537

   PIN n_125551
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 25.01 0.163 25.038 ;
      END
   END n_125551

   PIN n_12570
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 85.618 0.163 85.646 ;
      END
   END n_12570

   PIN n_125714
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 168.626 122.077 168.654 122.24 ;
      END
   END n_125714

   PIN n_125785
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.626 122.077 80.654 122.24 ;
      END
   END n_125785

   PIN n_126191
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.106 122.077 85.134 122.24 ;
      END
   END n_126191

   PIN n_126306
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 313.23 114.61 313.394 114.638 ;
      END
   END n_126306

   PIN n_126307
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 113.33 313.394 113.358 ;
      END
   END n_126307

   PIN n_126587
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.442 122.077 11.47 122.24 ;
      END
   END n_126587

   PIN n_126600
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.242 122.077 80.27 122.24 ;
      END
   END n_126600

   PIN n_126601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.778 122.077 81.806 122.24 ;
      END
   END n_126601

   PIN n_12712
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 141.746 122.077 141.774 122.24 ;
      END
   END n_12712

   PIN n_127297
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.426 0.163 117.454 ;
      END
   END n_127297

   PIN n_127737
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.106 122.077 245.134 122.24 ;
      END
   END n_127737

   PIN n_127742
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 237.682 122.077 237.71 122.24 ;
      END
   END n_127742

   PIN n_127891
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.234 0.163 117.262 ;
      END
   END n_127891

   PIN n_128372
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.49 0.163 117.518 ;
      END
   END n_128372

   PIN n_128584
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 245.554 122.077 245.582 122.24 ;
      END
   END n_128584

   PIN n_128848
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 303.218 122.077 303.246 122.24 ;
      END
   END n_128848

   PIN n_128849
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 312.114 122.077 312.142 122.24 ;
      END
   END n_128849

   PIN n_128989
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.074 122.077 65.102 122.24 ;
      END
   END n_128989

   PIN n_129129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.114 0.163 48.142 ;
      END
   END n_129129

   PIN n_129403
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.874 0.163 117.902 ;
      END
   END n_129403

   PIN n_129491
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 312.178 122.077 312.206 122.24 ;
      END
   END n_129491

   PIN n_129545
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.762 122.077 3.79 122.24 ;
      END
   END n_129545

   PIN n_129619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 264.882 122.077 264.91 122.24 ;
      END
   END n_129619

   PIN n_129824
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.522 0.163 105.55 ;
      END
   END n_129824

   PIN n_129826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 117.17 0.163 117.198 ;
      END
   END n_129826

   PIN n_129827
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 312.242 122.077 312.27 122.24 ;
      END
   END n_129827

   PIN n_129828
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.01 122.077 65.038 122.24 ;
      END
   END n_129828

   PIN n_129897
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.826 122.077 3.854 122.24 ;
      END
   END n_129897

   PIN n_130137
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 60.978 313.394 61.006 ;
      END
   END n_130137

   PIN n_130202
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 28.978 313.394 29.006 ;
      END
   END n_130202

   PIN n_130204
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 117.17 313.394 117.198 ;
      END
   END n_130204

   PIN n_130594
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 141.81 122.077 141.838 122.24 ;
      END
   END n_130594

   PIN n_130626
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 287.858 122.077 287.886 122.24 ;
      END
   END n_130626

   PIN n_131059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 284.082 122.077 284.11 122.24 ;
      END
   END n_131059

   PIN n_131060
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 260.978 122.077 261.006 122.24 ;
      END
   END n_131060

   PIN n_131305
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.226 0.163 98.254 ;
      END
   END n_131305

   PIN n_131421
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 287.922 122.077 287.95 122.24 ;
      END
   END n_131421

   PIN n_131475
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.738 0.163 82.766 ;
      END
   END n_131475

   PIN n_132026
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.834 122.077 110.862 122.24 ;
      END
   END n_132026

   PIN n_132027
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.89 122.077 115.918 122.24 ;
      END
   END n_132027

   PIN n_132085
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.65 122.077 145.678 122.24 ;
      END
   END n_132085

   PIN n_132293
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.538 122.077 7.566 122.24 ;
      END
   END n_132293

   PIN n_132825
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.25 122.077 107.278 122.24 ;
      END
   END n_132825

   PIN n_132870
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 197.874 122.077 197.902 122.24 ;
      END
   END n_132870

   PIN n_133002
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.97 0.163 113.998 ;
      END
   END n_133002

   PIN n_133183
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 105.842 0.163 105.87 ;
      END
   END n_133183

   PIN n_133738
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 90.29 0.163 90.318 ;
      END
   END n_133738

   PIN n_133859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 312.178 122.077 312.206 122.24 ;
      END
   END n_133859

   PIN n_133940
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 312.306 122.077 312.334 122.24 ;
      END
   END n_133940

   PIN n_134182
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 115.506 122.077 115.534 122.24 ;
      END
   END n_134182

   PIN n_134553
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 306.994 122.077 307.022 122.24 ;
      END
   END n_134553

   PIN n_134648
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 312.37 122.077 312.398 122.24 ;
      END
   END n_134648

   PIN n_134804
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.346 122.077 111.374 122.24 ;
      END
   END n_134804

   PIN n_135056
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.714 0.163 113.742 ;
      END
   END n_135056

   PIN n_135073
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.514 0.163 78.542 ;
      END
   END n_135073

   PIN n_135074
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.578 0.163 78.606 ;
      END
   END n_135074

   PIN n_135796
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 299.314 122.077 299.342 122.24 ;
      END
   END n_135796

   PIN n_135808
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 173.17 122.077 173.198 122.24 ;
      END
   END n_135808

   PIN n_136154
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 280.242 122.077 280.27 122.24 ;
      END
   END n_136154

   PIN n_136201
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.138 122.077 57.166 122.24 ;
      END
   END n_136201

   PIN n_136203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.338 122.077 60.366 122.24 ;
      END
   END n_136203

   PIN n_136211
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.266 122.077 57.294 122.24 ;
      END
   END n_136211

   PIN n_136212
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.33 122.077 57.358 122.24 ;
      END
   END n_136212

   PIN n_136268
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 134.13 122.077 134.158 122.24 ;
      END
   END n_136268

   PIN n_136598
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 284.146 122.077 284.174 122.24 ;
      END
   END n_136598

   PIN n_136630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 276.274 122.077 276.302 122.24 ;
      END
   END n_136630

   PIN n_136660
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.394 0.163 17.422 ;
      END
   END n_136660

   PIN n_136842
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.266 0.163 17.294 ;
      END
   END n_136842

   PIN n_136875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.482 122.077 186.51 122.24 ;
      END
   END n_136875

   PIN n_136876
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 179.058 122.077 179.086 122.24 ;
      END
   END n_136876

   PIN n_136887
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.21 122.077 180.238 122.24 ;
      END
   END n_136887

   PIN n_137597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 264.69 122.077 264.718 122.24 ;
      END
   END n_137597

   PIN n_14162
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 128.178 122.077 128.206 122.24 ;
      END
   END n_14162

   PIN n_143063
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 117.554 0.163 117.582 ;
      END
   END n_143063

   PIN n_143692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.418 122.077 130.446 122.24 ;
      END
   END n_143692

   PIN n_143725
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.258 0.163 86.286 ;
      END
   END n_143725

   PIN n_143810
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 153.394 122.077 153.422 122.24 ;
      END
   END n_143810

   PIN n_143811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.21 122.077 220.238 122.24 ;
      END
   END n_143811

   PIN n_14682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.29 0.163 98.318 ;
      END
   END n_14682

   PIN n_16033
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 168.754 122.077 168.782 122.24 ;
      END
   END n_16033

   PIN n_16164
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 114.93 122.077 114.958 122.24 ;
      END
   END n_16164

   PIN n_16207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 122.674 122.077 122.702 122.24 ;
      END
   END n_16207

   PIN n_16296
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 214.706 122.077 214.734 122.24 ;
      END
   END n_16296

   PIN n_18629
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.714 122.077 241.742 122.24 ;
      END
   END n_18629

   PIN n_18630
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.266 122.077 241.294 122.24 ;
      END
   END n_18630

   PIN n_18732
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 214.834 122.077 214.862 122.24 ;
      END
   END n_18732

   PIN n_18908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.194 122.077 38.222 122.24 ;
      END
   END n_18908

   PIN n_18997
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 168.69 122.077 168.718 122.24 ;
      END
   END n_18997

   PIN n_19022
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.65 122.077 241.678 122.24 ;
      END
   END n_19022

   PIN n_19642
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.73 122.077 7.758 122.24 ;
      END
   END n_19642

   PIN n_20025
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 122.738 122.077 122.766 122.24 ;
      END
   END n_20025

   PIN n_20054
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.874 0.163 109.902 ;
      END
   END n_20054

   PIN n_20260
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.026 122.077 207.054 122.24 ;
      END
   END n_20260

   PIN n_20282
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.13 122.077 134.158 122.24 ;
      END
   END n_20282

   PIN n_20329
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.178 122.077 224.206 122.24 ;
      END
   END n_20329

   PIN n_20334
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 183.986 122.077 184.014 122.24 ;
      END
   END n_20334

   PIN n_20442
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.186 122.077 203.214 122.24 ;
      END
   END n_20442

   PIN n_20443
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.25 122.077 203.278 122.24 ;
      END
   END n_20443

   PIN n_20690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.314 122.077 203.342 122.24 ;
      END
   END n_20690

   PIN n_20855
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 284.082 122.077 284.11 122.24 ;
      END
   END n_20855

   PIN n_20865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 230.066 122.077 230.094 122.24 ;
      END
   END n_20865

   PIN n_20867
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 137.842 122.077 137.87 122.24 ;
      END
   END n_20867

   PIN n_20880
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 130.29 122.077 130.318 122.24 ;
      END
   END n_20880

   PIN n_21104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 185.202 122.077 185.23 122.24 ;
      END
   END n_21104

   PIN n_21252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 184.242 122.077 184.27 122.24 ;
      END
   END n_21252

   PIN n_21408
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 210.994 122.077 211.022 122.24 ;
      END
   END n_21408

   PIN n_21512
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.506 122.077 67.534 122.24 ;
      END
   END n_21512

   PIN n_21514
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.762 122.077 67.79 122.24 ;
      END
   END n_21514

   PIN n_21917
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 313.23 117.682 313.394 117.71 ;
      END
   END n_21917

   PIN n_22013
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 210.866 122.077 210.894 122.24 ;
      END
   END n_22013

   PIN n_22014
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 210.93 122.077 210.958 122.24 ;
      END
   END n_22014

   PIN n_22238
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.41 122.077 79.438 122.24 ;
      END
   END n_22238

   PIN n_22308
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.09 122.077 207.118 122.24 ;
      END
   END n_22308

   PIN n_22322
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.218 122.077 207.246 122.24 ;
      END
   END n_22322

   PIN n_22555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.57 122.077 195.598 122.24 ;
      END
   END n_22555

   PIN n_22556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 198.706 122.077 198.734 122.24 ;
      END
   END n_22556

   PIN n_22569
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 184.178 122.077 184.206 122.24 ;
      END
   END n_22569

   PIN n_22576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 184.05 122.077 184.078 122.24 ;
      END
   END n_22576

   PIN n_23134
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.746 122.077 229.774 122.24 ;
      END
   END n_23134

   PIN n_23144
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 222.386 122.077 222.414 122.24 ;
      END
   END n_23144

   PIN n_23481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 199.794 122.077 199.822 122.24 ;
      END
   END n_23481

   PIN n_23793
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 141.874 122.077 141.902 122.24 ;
      END
   END n_23793

   PIN n_23795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 141.874 122.077 141.902 122.24 ;
      END
   END n_23795

   PIN n_24123
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 205.426 122.077 205.454 122.24 ;
      END
   END n_24123

   PIN n_24149
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 221.298 122.077 221.326 122.24 ;
      END
   END n_24149

   PIN n_24687
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.826 122.077 195.854 122.24 ;
      END
   END n_24687

   PIN n_24724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 161.01 122.077 161.038 122.24 ;
      END
   END n_24724

   PIN n_24767
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 222.514 122.077 222.542 122.24 ;
      END
   END n_24767

   PIN n_24775
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 248.498 122.077 248.526 122.24 ;
      END
   END n_24775

   PIN n_24776
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.594 122.077 220.622 122.24 ;
      END
   END n_24776

   PIN n_24781
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 164.85 122.077 164.878 122.24 ;
      END
   END n_24781

   PIN n_25313
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 220.53 122.077 220.558 122.24 ;
      END
   END n_25313

   PIN n_25456
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.954 122.077 3.982 122.24 ;
      END
   END n_25456

   PIN n_26039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 191.794 122.077 191.822 122.24 ;
      END
   END n_26039

   PIN n_26051
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 139.378 122.077 139.406 122.24 ;
      END
   END n_26051

   PIN n_27859
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 109.49 313.394 109.518 ;
      END
   END n_27859

   PIN n_3190
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.938 0.163 109.966 ;
      END
   END n_3190

   PIN n_32795
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.034 122.077 42.062 122.24 ;
      END
   END n_32795

   PIN n_33263
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 303.09 122.077 303.118 122.24 ;
      END
   END n_33263

   PIN n_3333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 117.234 0.163 117.262 ;
      END
   END n_3333

   PIN n_33852
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.45 122.077 126.478 122.24 ;
      END
   END n_33852

   PIN n_34115
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 102.13 0.163 102.158 ;
      END
   END n_34115

   PIN n_34197
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.578 122.077 86.606 122.24 ;
      END
   END n_34197

   PIN n_34198
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 84.21 122.077 84.238 122.24 ;
      END
   END n_34198

   PIN n_34301
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.322 0.163 86.35 ;
      END
   END n_34301

   PIN n_34458
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 312.562 122.077 312.59 122.24 ;
      END
   END n_34458

   PIN n_34462
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.906 0.163 105.934 ;
      END
   END n_34462

   PIN n_34463
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.546 0.163 98.574 ;
      END
   END n_34463

   PIN n_34772
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.466 122.077 60.494 122.24 ;
      END
   END n_34772

   PIN n_34826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 235.378 122.077 235.406 122.24 ;
      END
   END n_34826

   PIN n_34941
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.354 0.163 98.382 ;
      END
   END n_34941

   PIN n_35030
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.514 122.077 30.542 122.24 ;
      END
   END n_35030

   PIN n_35071
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 303.154 122.077 303.182 122.24 ;
      END
   END n_35071

   PIN n_36024
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 307.122 122.077 307.15 122.24 ;
      END
   END n_36024

   PIN n_3760
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.354 0.163 90.382 ;
      END
   END n_3760

   PIN n_5402
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 181.554 122.077 181.582 122.24 ;
      END
   END n_5402

   PIN n_5571
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 161.074 122.077 161.102 122.24 ;
      END
   END n_5571

   PIN n_7597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.586 122.077 241.614 122.24 ;
      END
   END n_7597

   PIN n_7782
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 83.442 0.163 83.47 ;
      END
   END n_7782

   PIN n_7815
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.89 122.077 3.918 122.24 ;
      END
   END n_7815

   PIN n_7857
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.042 0.163 45.07 ;
      END
   END n_7857

   PIN n_9933
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 218.61 122.077 218.638 122.24 ;
      END
   END n_9933

   PIN FE_OCPN19344_n_142919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.154 122.077 207.182 122.24 ;
      END
   END FE_OCPN19344_n_142919

   PIN FE_OFN10229_b_2_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 85.298 0.163 85.326 ;
      END
   END FE_OFN10229_b_2_6_2

   PIN FE_OFN10255_b_2_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.682 122.077 93.71 122.24 ;
      END
   END FE_OFN10255_b_2_4_7

   PIN FE_OFN10258_b_2_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 117.682 0.163 117.71 ;
      END
   END FE_OFN10258_b_2_4_5

   PIN FE_OFN10270_b_2_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.194 0.163 94.222 ;
      END
   END FE_OFN10270_b_2_4_1

   PIN FE_OFN10273_b_2_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.506 122.077 11.534 122.24 ;
      END
   END FE_OFN10273_b_2_4_0

   PIN FE_OFN10291_b_2_2_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.018 122.077 36.046 122.24 ;
      END
   END FE_OFN10291_b_2_2_4

   PIN FE_OFN1088_n_20334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 187.89 122.077 187.918 122.24 ;
      END
   END FE_OFN1088_n_20334

   PIN FE_OFN1106_n_19671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 209.522 122.077 209.55 122.24 ;
      END
   END FE_OFN1106_n_19671

   PIN FE_OFN11336_n_143645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.226 0.163 90.254 ;
      END
   END FE_OFN11336_n_143645

   PIN FE_OFN11351_n_140257
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 117.49 0.163 117.518 ;
      END
   END FE_OFN11351_n_140257

   PIN FE_OFN11361_n_143059
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 143.218 122.077 143.246 122.24 ;
      END
   END FE_OFN11361_n_143059

   PIN FE_OFN11368_n_143045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 175.73 122.077 175.758 122.24 ;
      END
   END FE_OFN11368_n_143045

   PIN FE_OFN11370_n_143045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.258 122.077 134.286 122.24 ;
      END
   END FE_OFN11370_n_143045

   PIN FE_OFN11397_n_140245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.674 0.163 90.702 ;
      END
   END FE_OFN11397_n_140245

   PIN FE_OFN11427_n_142905
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.066 122.077 166.094 122.24 ;
      END
   END FE_OFN11427_n_142905

   PIN FE_OFN11432_n_142919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.442 122.077 211.47 122.24 ;
      END
   END FE_OFN11432_n_142919

   PIN FE_OFN11590_n_143231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.602 122.077 7.63 122.24 ;
      END
   END FE_OFN11590_n_143231

   PIN FE_OFN11596_n_112428
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.81 0.163 93.838 ;
      END
   END FE_OFN11596_n_112428

   PIN FE_OFN11705_n_142947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.642 0.163 118.67 ;
      END
   END FE_OFN11705_n_142947

   PIN FE_OFN11865_n_143230
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.106 0.163 61.134 ;
      END
   END FE_OFN11865_n_143230

   PIN FE_OFN11869_n_143229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 75.058 0.163 75.086 ;
      END
   END FE_OFN11869_n_143229

   PIN FE_OFN11871_n_143229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 107.378 122.077 107.406 122.24 ;
      END
   END FE_OFN11871_n_143229

   PIN FE_OFN11875_n_143227
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.098 122.077 138.126 122.24 ;
      END
   END FE_OFN11875_n_143227

   PIN FE_OFN11889_n_143104
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.522 0.163 97.55 ;
      END
   END FE_OFN11889_n_143104

   PIN FE_OFN11896_n_143102
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.178 122.077 88.206 122.24 ;
      END
   END FE_OFN11896_n_143102

   PIN FE_OFN11917_n_143048
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.322 0.163 118.35 ;
      END
   END FE_OFN11917_n_143048

   PIN FE_OFN12298_n_111727
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 139.314 122.077 139.342 122.24 ;
      END
   END FE_OFN12298_n_111727

   PIN FE_OFN12309_n_111875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.978 122.158 101.006 122.24 ;
      END
   END FE_OFN12309_n_111875

   PIN FE_OFN12318_n_111878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.13 0.163 94.158 ;
      END
   END FE_OFN12318_n_111878

   PIN FE_OFN12322_n_112427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 105.714 0.163 105.742 ;
      END
   END FE_OFN12322_n_112427

   PIN FE_OFN12325_n_112470
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.666 122.077 7.694 122.24 ;
      END
   END FE_OFN12325_n_112470

   PIN FE_OFN12332_n_137473
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.93 122.077 18.958 122.24 ;
      END
   END FE_OFN12332_n_137473

   PIN FE_OFN12348_n_142991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 106.098 122.077 106.126 122.24 ;
      END
   END FE_OFN12348_n_142991

   PIN FE_OFN12350_n_142991
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 85.426 0.163 85.454 ;
      END
   END FE_OFN12350_n_142991

   PIN FE_OFN12378_n_142908
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.09 122.077 15.118 122.24 ;
      END
   END FE_OFN12378_n_142908

   PIN FE_OFN12597_n_111737
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 69.81 0.163 69.838 ;
      END
   END FE_OFN12597_n_111737

   PIN FE_OFN12599_n_111738
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.458 0.163 105.486 ;
      END
   END FE_OFN12599_n_111738

   PIN FE_OFN12609_n_112606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.002 0.082 94.03 ;
      END
   END FE_OFN12609_n_112606

   PIN FE_OFN12611_n_112608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.362 122.077 109.39 122.24 ;
      END
   END FE_OFN12611_n_112608

   PIN FE_OFN12616_n_112689
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 101.618 0.163 101.646 ;
      END
   END FE_OFN12616_n_112689

   PIN FE_OFN12621_n_112690
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.994 122.077 19.022 122.24 ;
      END
   END FE_OFN12621_n_112690

   PIN FE_OFN12627_n_143646
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.482 0.163 82.51 ;
      END
   END FE_OFN12627_n_143646

   PIN FE_OFN12655_n_111913
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 85.362 0.163 85.39 ;
      END
   END FE_OFN12655_n_111913

   PIN FE_OFN12715_n_142865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 264.754 122.077 264.782 122.24 ;
      END
   END FE_OFN12715_n_142865

   PIN FE_OFN12960_n_111998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 264.69 122.158 264.718 122.24 ;
      END
   END FE_OFN12960_n_111998

   PIN FE_OFN12965_n_112000
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 211.634 122.077 211.662 122.24 ;
      END
   END FE_OFN12965_n_112000

   PIN FE_OFN12970_n_112611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 218.738 122.158 218.766 122.24 ;
      END
   END FE_OFN12970_n_112611

   PIN FE_OFN12985_n_112681
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 287.73 122.077 287.758 122.24 ;
      END
   END FE_OFN12985_n_112681

   PIN FE_OFN13013_n_142950
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 114.738 0.163 114.766 ;
      END
   END FE_OFN13013_n_142950

   PIN FE_OFN13023_n_142949
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 78.77 0.163 78.798 ;
      END
   END FE_OFN13023_n_142949

   PIN FE_OFN13543_n_143609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 287.794 122.077 287.822 122.24 ;
      END
   END FE_OFN13543_n_143609

   PIN FE_OFN13547_n_112256
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.034 122.077 226.062 122.24 ;
      END
   END FE_OFN13547_n_112256

   PIN FE_OFN13556_n_143397
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.618 0.163 93.646 ;
      END
   END FE_OFN13556_n_143397

   PIN FE_OFN13659_n_112318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 272.434 122.077 272.462 122.24 ;
      END
   END FE_OFN13659_n_112318

   PIN FE_OFN13700_n_143384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 295.602 122.077 295.63 122.24 ;
      END
   END FE_OFN13700_n_143384

   PIN FE_OFN13708_n_143383
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 280.178 122.077 280.206 122.24 ;
      END
   END FE_OFN13708_n_143383

   PIN FE_OFN13818_n_112257
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 284.018 122.077 284.046 122.24 ;
      END
   END FE_OFN13818_n_112257

   PIN FE_OFN14269_n_140244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.258 0.163 118.286 ;
      END
   END FE_OFN14269_n_140244

   PIN FE_OFN14270_n_140244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.61 0.163 90.638 ;
      END
   END FE_OFN14270_n_140244

   PIN FE_OFN15080_n_19611
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 148.594 122.077 148.622 122.24 ;
      END
   END FE_OFN15080_n_19611

   PIN FE_OFN15155_n_23384
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.73 122.077 207.758 122.24 ;
      END
   END FE_OFN15155_n_23384

   PIN FE_OFN15251_n_39084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.922 122.077 311.95 122.24 ;
      END
   END FE_OFN15251_n_39084

   PIN FE_OFN16362_b_2_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.162 0.163 90.19 ;
      END
   END FE_OFN16362_b_2_6_1

   PIN FE_OFN16770_n_16098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.002 122.077 238.03 122.24 ;
      END
   END FE_OFN16770_n_16098

   PIN FE_OFN16941_n_135332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 207.09 122.077 207.118 122.24 ;
      END
   END FE_OFN16941_n_135332

   PIN FE_OFN17141_n_22815
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.314 0.163 67.342 ;
      END
   END FE_OFN17141_n_22815

   PIN FE_OFN17145_n_22232
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.41 0.163 63.438 ;
      END
   END FE_OFN17145_n_22232

   PIN FE_OFN17169_n_16270
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.458 0.163 97.486 ;
      END
   END FE_OFN17169_n_16270

   PIN FE_OFN17207_n_21410
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.25 0.163 67.278 ;
      END
   END FE_OFN17207_n_21410

   PIN FE_OFN17264_n_140245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 295.538 122.077 295.566 122.24 ;
      END
   END FE_OFN17264_n_140245

   PIN FE_OFN18602_b_2_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 94.066 0.163 94.094 ;
      END
   END FE_OFN18602_b_2_6_0

   PIN FE_OFN18750_n_112550
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.226 122.077 130.254 122.24 ;
      END
   END FE_OFN18750_n_112550

   PIN FE_OFN18809_n_143645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.722 122.077 212.75 122.24 ;
      END
   END FE_OFN18809_n_143645

   PIN FE_OFN19061_n_21194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.266 122.077 73.294 122.24 ;
      END
   END FE_OFN19061_n_21194

   PIN FE_OFN2152_n_19668
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.906 122.077 145.934 122.24 ;
      END
   END FE_OFN2152_n_19668

   PIN FE_OFN2159_n_19626
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.386 122.077 126.414 122.24 ;
      END
   END FE_OFN2159_n_19626

   PIN FE_OFN2284_n_19629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.762 122.077 91.79 122.24 ;
      END
   END FE_OFN2284_n_19629

   PIN FE_OFN3204_n_14458
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 187.634 122.077 187.662 122.24 ;
      END
   END FE_OFN3204_n_14458

   PIN FE_OFN3244_n_19948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.114 122.077 88.142 122.24 ;
      END
   END FE_OFN3244_n_19948

   PIN FE_OFN3293_n_8246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.866 0.163 74.894 ;
      END
   END FE_OFN3293_n_8246

   PIN FE_OFN3382_n_14610
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.65 0.163 97.678 ;
      END
   END FE_OFN3382_n_14610

   PIN FE_OFN3441_n_12341
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.026 0.163 71.054 ;
      END
   END FE_OFN3441_n_12341

   PIN FE_OFN3505_n_12951
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.05 0.163 48.078 ;
      END
   END FE_OFN3505_n_12951

   PIN FE_OFN3587_n_142906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.81 122.077 45.838 122.24 ;
      END
   END FE_OFN3587_n_142906

   PIN FE_OFN3683_n_142948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.578 0.163 94.606 ;
      END
   END FE_OFN3683_n_142948

   PIN FE_OFN3701_n_143060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.618 0.163 77.646 ;
      END
   END FE_OFN3701_n_143060

   PIN FE_OFN3720_n_143241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 121.906 122.077 121.934 122.24 ;
      END
   END FE_OFN3720_n_143241

   PIN FE_OFN3726_n_143241
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 89.906 0.163 89.934 ;
      END
   END FE_OFN3726_n_143241

   PIN FE_OFN3737_n_143396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.746 0.163 101.774 ;
      END
   END FE_OFN3737_n_143396

   PIN FE_OFN3743_n_143551
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.354 0.163 82.382 ;
      END
   END FE_OFN3743_n_143551

   PIN FE_OFN3751_n_143549
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.298 0.163 101.326 ;
      END
   END FE_OFN3751_n_143549

   PIN FE_OFN596_n_8407
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 199.41 122.077 199.438 122.24 ;
      END
   END FE_OFN596_n_8407

   PIN FE_OFN700_n_22202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 153.202 122.077 153.23 122.24 ;
      END
   END FE_OFN700_n_22202

   PIN FE_OFN791_n_19612
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.426 122.077 245.454 122.24 ;
      END
   END FE_OFN791_n_19612

   PIN FE_OFN794_n_20260
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 210.802 122.077 210.83 122.24 ;
      END
   END FE_OFN794_n_20260

   PIN FE_OFN832_n_22177
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 203.314 122.077 203.342 122.24 ;
      END
   END FE_OFN832_n_22177

   PIN FE_OFN9231_delay_add_ln34_unr2_unr3_stage2_stallmux_q_15_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 167.346 122.077 167.374 122.24 ;
      END
   END FE_OFN9231_delay_add_ln34_unr2_unr3_stage2_stallmux_q_15_

   PIN add_5900_51_n_88
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 260.978 122.077 261.006 122.24 ;
      END
   END add_5900_51_n_88

   PIN b_0_2_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.312 46.258 313.394 46.286 ;
      END
   END b_0_2_0

   PIN b_0_2_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 214.386 122.158 214.414 122.24 ;
      END
   END b_0_2_1

   PIN b_0_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.312 31.282 313.394 31.31 ;
      END
   END b_0_2_2

   PIN b_0_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.312 19.89 313.394 19.918 ;
      END
   END b_0_2_3

   PIN b_0_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 222.706 122.158 222.734 122.24 ;
      END
   END b_0_4_1

   PIN b_0_6_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.312 40.05 313.394 40.078 ;
      END
   END b_0_6_0

   PIN b_0_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 222.578 122.158 222.606 122.24 ;
      END
   END b_0_6_1

   PIN b_0_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.312 12.658 313.394 12.686 ;
      END
   END b_0_6_2

   PIN b_0_6_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 28.658 313.394 28.686 ;
      END
   END b_0_6_5

   PIN b_1_9_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 241.842 122.158 241.87 122.24 ;
      END
   END b_1_9_0

   PIN b_2_2_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.21 0.0 92.238 0.163 ;
      END
   END b_2_2_0

   PIN b_2_2_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 110.066 0.163 110.094 ;
      END
   END b_2_2_1

   PIN b_2_2_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.49 0.0 45.518 0.163 ;
      END
   END b_2_2_11

   PIN b_2_2_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 115.122 0.0 115.15 0.163 ;
      END
   END b_2_2_2

   PIN b_2_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 112.562 0.0 112.59 0.163 ;
      END
   END b_2_2_3

   PIN b_2_2_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 110.258 0.163 110.286 ;
      END
   END b_2_2_4

   PIN b_2_2_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 108.978 0.163 109.006 ;
      END
   END b_2_2_5

   PIN b_2_2_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.13 0.163 102.158 ;
      END
   END b_2_2_6

   PIN b_2_2_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 106.034 0.163 106.062 ;
      END
   END b_2_2_7

   PIN b_2_2_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.386 0.163 118.414 ;
      END
   END b_2_2_8

   PIN b_2_4_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.778 122.077 145.806 122.24 ;
      END
   END b_2_4_0

   PIN b_2_4_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 85.426 0.163 85.454 ;
      END
   END b_2_4_1

   PIN b_2_4_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 141.362 122.077 141.39 122.24 ;
      END
   END b_2_4_11

   PIN b_2_4_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 110.002 0.163 110.03 ;
      END
   END b_2_4_12

   PIN b_2_4_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 108.658 0.0 108.686 0.163 ;
      END
   END b_2_4_13

   PIN b_2_4_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.554 0.0 69.582 0.163 ;
      END
   END b_2_4_2

   PIN b_2_4_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 144.562 122.077 144.59 122.24 ;
      END
   END b_2_4_3

   PIN b_2_4_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.25 122.077 139.278 122.24 ;
      END
   END b_2_4_4

   PIN b_2_4_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.794 0.0 87.822 0.163 ;
      END
   END b_2_4_5

   PIN b_2_4_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 94.77 0.0 94.798 0.163 ;
      END
   END b_2_4_6

   PIN b_2_4_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.21 122.077 124.238 122.24 ;
      END
   END b_2_4_7

   PIN b_2_4_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 102.002 0.163 102.03 ;
      END
   END b_2_4_8

   PIN b_2_6_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 136.434 122.077 136.462 122.24 ;
      END
   END b_2_6_1

   PIN b_2_6_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 138.162 122.077 138.19 122.24 ;
      END
   END b_2_6_10

   PIN b_2_6_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.69 122.077 120.718 122.24 ;
      END
   END b_2_6_11

   PIN b_2_6_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 130.354 122.077 130.382 122.24 ;
      END
   END b_2_6_12

   PIN b_2_6_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.258 0.163 94.286 ;
      END
   END b_2_6_13

   PIN b_2_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 132.978 122.077 133.006 122.24 ;
      END
   END b_2_6_2

   PIN b_2_6_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.882 122.077 152.91 122.24 ;
      END
   END b_2_6_3

   PIN b_2_6_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 154.098 122.077 154.126 122.24 ;
      END
   END b_2_6_4

   PIN b_2_6_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.37 122.077 160.398 122.24 ;
      END
   END b_2_6_7

   PIN b_2_6_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.002 0.0 126.03 0.163 ;
      END
   END b_2_6_9

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 205.106 122.158 205.134 122.24 ;
      END
   END ispd_clk

   PIN mul_4370_72_n_149
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.506 122.077 307.534 122.24 ;
      END
   END mul_4370_72_n_149

   PIN mul_4370_72_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 257.074 122.077 257.102 122.24 ;
      END
   END mul_4370_72_n_50

   PIN mul_4370_72_n_66
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.858 122.077 311.886 122.24 ;
      END
   END mul_4370_72_n_66

   PIN mul_4370_72_n_793
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 310.962 122.077 310.99 122.24 ;
      END
   END mul_4370_72_n_793

   PIN mul_4370_72_n_840
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.25 122.077 307.278 122.24 ;
      END
   END mul_4370_72_n_840

   PIN mul_4377_72_n_106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 248.434 122.077 248.462 122.24 ;
      END
   END mul_4377_72_n_106

   PIN mul_4377_72_n_114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 149.618 122.077 149.646 122.24 ;
      END
   END mul_4377_72_n_114

   PIN mul_4377_72_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 230.194 122.077 230.222 122.24 ;
      END
   END mul_4377_72_n_116

   PIN mul_4665_72_n_244
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.266 0.163 113.294 ;
      END
   END mul_4665_72_n_244

   PIN mul_4665_72_n_330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.17 0.163 117.198 ;
      END
   END mul_4665_72_n_330

   PIN mul_4665_72_n_338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.082 0.163 44.11 ;
      END
   END mul_4665_72_n_338

   PIN mul_4665_72_n_339
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.306 0.163 40.334 ;
      END
   END mul_4665_72_n_339

   PIN mul_4667_72_n_334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 101.746 122.077 101.774 122.24 ;
      END
   END mul_4667_72_n_334

   PIN mul_4667_72_n_340
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 74.866 0.163 74.894 ;
      END
   END mul_4667_72_n_340

   PIN mul_4669_72_n_315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 101.938 0.163 101.966 ;
      END
   END mul_4669_72_n_315

   PIN mul_4669_72_n_340
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.282 0.163 63.31 ;
      END
   END mul_4669_72_n_340

   PIN mul_ln34_unr2_unr2_z_11_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.33 0.163 97.358 ;
      END
   END mul_ln34_unr2_unr2_z_11_

   PIN mul_ln34_unr2_unr5_z_13_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 61.042 0.163 61.07 ;
      END
   END mul_ln34_unr2_unr5_z_13_

   PIN mul_ln34_unr2_unr5_z_14_
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.106 0.163 45.134 ;
      END
   END mul_ln34_unr2_unr5_z_14_

   PIN n_10106
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.746 0.163 117.774 ;
      END
   END n_10106

   PIN n_10396
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.09 122.077 111.118 122.24 ;
      END
   END n_10396

   PIN n_10648
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.17 122.077 157.198 122.24 ;
      END
   END n_10648

   PIN n_10996
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 122.61 122.077 122.638 122.24 ;
      END
   END n_10996

   PIN n_10998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 264.626 122.077 264.654 122.24 ;
      END
   END n_10998

   PIN n_111930
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 223.858 122.077 223.886 122.24 ;
      END
   END n_111930

   PIN n_112180
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.314 122.077 11.342 122.24 ;
      END
   END n_112180

   PIN n_112566
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.858 122.077 7.886 122.24 ;
      END
   END n_112566

   PIN n_112607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.218 122.158 15.246 122.24 ;
      END
   END n_112607

   PIN n_112707
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.794 122.077 311.822 122.24 ;
      END
   END n_112707

   PIN n_112826
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.25 122.077 11.278 122.24 ;
      END
   END n_112826

   PIN n_112827
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.186 122.077 11.214 122.24 ;
      END
   END n_112827

   PIN n_112875
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.218 122.077 15.246 122.24 ;
      END
   END n_112875

   PIN n_112887
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 283.954 122.077 283.982 122.24 ;
      END
   END n_112887

   PIN n_112910
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 312.306 122.077 312.334 122.24 ;
      END
   END n_112910

   PIN n_112911
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 310.898 122.077 310.926 122.24 ;
      END
   END n_112911

   PIN n_112930
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 226.226 122.077 226.254 122.24 ;
      END
   END n_112930

   PIN n_113050
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 295.346 122.077 295.374 122.24 ;
      END
   END n_113050

   PIN n_113218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 114.674 0.163 114.702 ;
      END
   END n_113218

   PIN n_113364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 54.578 313.394 54.606 ;
      END
   END n_113364

   PIN n_113365
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 117.106 313.394 117.134 ;
      END
   END n_113365

   PIN n_113366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 191.218 122.077 191.246 122.24 ;
      END
   END n_113366

   PIN n_113426
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 295.538 122.077 295.566 122.24 ;
      END
   END n_113426

   PIN n_113502
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.634 122.077 3.662 122.24 ;
      END
   END n_113502

   PIN n_113544
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.578 0.163 118.606 ;
      END
   END n_113544

   PIN n_113546
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.458 0.163 113.486 ;
      END
   END n_113546

   PIN n_113561
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.098 0.163 98.126 ;
      END
   END n_113561

   PIN n_113602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 313.23 105.65 313.394 105.678 ;
      END
   END n_113602

   PIN n_113603
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 53.298 313.394 53.326 ;
      END
   END n_113603

   PIN n_113699
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 93.938 0.163 93.966 ;
      END
   END n_113699

   PIN n_113855
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.474 122.077 7.502 122.24 ;
      END
   END n_113855

   PIN n_113856
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 93.874 0.163 93.902 ;
      END
   END n_113856

   PIN n_113866
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 90.098 0.163 90.126 ;
      END
   END n_113866

   PIN n_113926
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.29 0.163 82.318 ;
      END
   END n_113926

   PIN n_113994
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.162 0.163 114.19 ;
      END
   END n_113994

   PIN n_114084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.802 0.163 74.83 ;
      END
   END n_114084

   PIN n_114198
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.122 0.163 67.15 ;
      END
   END n_114198

   PIN n_114263
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.834 0.163 78.862 ;
      END
   END n_114263

   PIN n_114274
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.682 0.163 117.71 ;
      END
   END n_114274

   PIN n_114292
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 295.282 122.077 295.31 122.24 ;
      END
   END n_114292

   PIN n_114416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.386 0.163 86.414 ;
      END
   END n_114416

   PIN n_114432
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.034 0.163 98.062 ;
      END
   END n_114432

   PIN n_114581
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 292.914 122.077 292.942 122.24 ;
      END
   END n_114581

   PIN n_114701
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.394 0.163 105.422 ;
      END
   END n_114701

   PIN n_115305
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.106 0.163 117.134 ;
      END
   END n_115305

   PIN n_11535
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.026 122.077 111.054 122.24 ;
      END
   END n_11535

   PIN n_115461
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.298 0.163 53.326 ;
      END
   END n_115461

   PIN n_115480
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 47.986 0.163 48.014 ;
      END
   END n_115480

   PIN n_115635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.538 122.077 7.566 122.24 ;
      END
   END n_115635

   PIN n_115636
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.77 122.077 22.798 122.24 ;
      END
   END n_115636

   PIN n_116469
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.474 122.077 7.502 122.24 ;
      END
   END n_116469

   PIN n_117228
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.842 122.077 145.87 122.24 ;
      END
   END n_117228

   PIN n_117236
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 244.402 122.077 244.43 122.24 ;
      END
   END n_117236

   PIN n_117237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.73 122.077 311.758 122.24 ;
      END
   END n_117237

   PIN n_117368
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 120.178 122.077 120.206 122.24 ;
      END
   END n_117368

   PIN n_117402
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 214.706 122.077 214.734 122.24 ;
      END
   END n_117402

   PIN n_117521
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.122 122.077 11.15 122.24 ;
      END
   END n_117521

   PIN n_118323
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.098 0.163 90.126 ;
      END
   END n_118323

   PIN n_119297
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.442 122.077 91.47 122.24 ;
      END
   END n_119297

   PIN n_119298
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.25 122.077 91.278 122.24 ;
      END
   END n_119298

   PIN n_119316
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.058 122.077 11.086 122.24 ;
      END
   END n_119316

   PIN n_119738
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.346 0.163 63.374 ;
      END
   END n_119738

   PIN n_119899
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.522 122.077 145.55 122.24 ;
      END
   END n_119899

   PIN n_119933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 313.23 117.106 313.394 117.134 ;
      END
   END n_119933

   PIN n_119934
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 53.362 313.394 53.39 ;
      END
   END n_119934

   PIN n_119959
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 249.33 122.077 249.358 122.24 ;
      END
   END n_119959

   PIN n_119983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 74.738 0.163 74.766 ;
      END
   END n_119983

   PIN n_120078
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.17 122.077 61.198 122.24 ;
      END
   END n_120078

   PIN n_120079
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.106 122.077 61.134 122.24 ;
      END
   END n_120079

   PIN n_120193
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 97.97 313.394 97.998 ;
      END
   END n_120193

   PIN n_120437
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 153.266 122.077 153.294 122.24 ;
      END
   END n_120437

   PIN n_120635
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.33 0.163 105.358 ;
      END
   END n_120635

   PIN n_120746
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 90.162 0.163 90.19 ;
      END
   END n_120746

   PIN n_120996
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.618 0.163 117.646 ;
      END
   END n_120996

   PIN n_121285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.666 122.077 311.694 122.24 ;
      END
   END n_121285

   PIN n_121633
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 246.834 122.077 246.862 122.24 ;
      END
   END n_121633

   PIN n_121772
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.866 122.077 82.894 122.24 ;
      END
   END n_121772

   PIN n_121803
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 313.23 94.13 313.394 94.158 ;
      END
   END n_121803

   PIN n_121832
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 291.698 122.077 291.726 122.24 ;
      END
   END n_121832

   PIN n_121834
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 272.37 122.077 272.398 122.24 ;
      END
   END n_121834

   PIN n_121906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.658 0.163 36.686 ;
      END
   END n_121906

   PIN n_121932
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 268.594 122.077 268.622 122.24 ;
      END
   END n_121932

   PIN n_121933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.738 122.077 242.766 122.24 ;
      END
   END n_121933

   PIN n_122107
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.842 0.163 97.87 ;
      END
   END n_122107

   PIN n_122555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 257.01 122.077 257.038 122.24 ;
      END
   END n_122555

   PIN n_122556
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 260.914 122.077 260.942 122.24 ;
      END
   END n_122556

   PIN n_12342
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.978 0.163 29.006 ;
      END
   END n_12342

   PIN n_123546
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 295.41 122.077 295.438 122.24 ;
      END
   END n_123546

   PIN n_123558
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 295.474 122.077 295.502 122.24 ;
      END
   END n_123558

   PIN n_123606
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.618 0.163 109.646 ;
      END
   END n_123606

   PIN n_123620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 268.53 122.077 268.558 122.24 ;
      END
   END n_123620

   PIN n_123678
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.514 122.077 62.542 122.24 ;
      END
   END n_123678

   PIN n_123759
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.442 122.077 307.47 122.24 ;
      END
   END n_123759

   PIN n_124048
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.546 0.163 90.574 ;
      END
   END n_124048

   PIN n_124617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.482 0.163 90.51 ;
      END
   END n_124617

   PIN n_124974
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.714 0.163 105.742 ;
      END
   END n_124974

   PIN n_124975
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.65 0.163 105.678 ;
      END
   END n_124975

   PIN n_125043
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 218.546 122.077 218.574 122.24 ;
      END
   END n_125043

   PIN n_125044
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 238.578 122.077 238.606 122.24 ;
      END
   END n_125044

   PIN n_125081
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.554 122.077 149.582 122.24 ;
      END
   END n_125081

   PIN n_125082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.49 122.077 149.518 122.24 ;
      END
   END n_125082

   PIN n_125769
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.602 122.077 311.63 122.24 ;
      END
   END n_125769

   PIN n_125781
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.282 122.077 311.31 122.24 ;
      END
   END n_125781

   PIN n_125786
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 312.242 122.077 312.27 122.24 ;
      END
   END n_125786

   PIN n_12587
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.77 0.163 78.798 ;
      END
   END n_12587

   PIN n_126291
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 69.298 313.394 69.326 ;
      END
   END n_126291

   PIN n_126292
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 74.93 313.394 74.958 ;
      END
   END n_126292

   PIN n_126559
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 109.426 313.394 109.454 ;
      END
   END n_126559

   PIN n_126560
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 20.658 313.394 20.686 ;
      END
   END n_126560

   PIN n_12711
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 177.778 122.077 177.806 122.24 ;
      END
   END n_12711

   PIN n_127736
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 245.17 122.077 245.198 122.24 ;
      END
   END n_127736

   PIN n_127873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 310.834 122.077 310.862 122.24 ;
      END
   END n_127873

   PIN n_127889
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.746 0.163 109.774 ;
      END
   END n_127889

   PIN n_127896
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 245.49 122.077 245.518 122.24 ;
      END
   END n_127896

   PIN n_127954
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.218 122.077 311.246 122.24 ;
      END
   END n_127954

   PIN n_128003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.45 0.163 94.478 ;
      END
   END n_128003

   PIN n_128515
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 257.01 122.077 257.038 122.24 ;
      END
   END n_128515

   PIN n_128527
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 235.25 122.077 235.278 122.24 ;
      END
   END n_128527

   PIN n_128971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.066 0.163 102.094 ;
      END
   END n_128971

   PIN n_128973
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 102.002 0.163 102.03 ;
      END
   END n_128973

   PIN n_129101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 89.842 0.163 89.87 ;
      END
   END n_129101

   PIN n_12956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 128.242 122.077 128.27 122.24 ;
      END
   END n_12956

   PIN n_130212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.874 0.163 93.902 ;
      END
   END n_130212

   PIN n_130734
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.586 0.163 97.614 ;
      END
   END n_130734

   PIN n_131017
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 76.978 0.163 77.006 ;
      END
   END n_131017

   PIN n_131069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 65.01 122.077 65.038 122.24 ;
      END
   END n_131069

   PIN n_131070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.074 122.077 65.102 122.24 ;
      END
   END n_131070

   PIN n_131430
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.722 0.163 20.75 ;
      END
   END n_131430

   PIN n_131641
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 72.754 122.077 72.782 122.24 ;
      END
   END n_131641

   PIN n_132252
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.642 122.077 110.67 122.24 ;
      END
   END n_132252

   PIN n_132417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.186 122.077 307.214 122.24 ;
      END
   END n_132417

   PIN n_132434
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.122 122.077 307.15 122.24 ;
      END
   END n_132434

   PIN n_132699
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.194 0.163 118.222 ;
      END
   END n_132699

   PIN n_132892
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.13 0.163 118.158 ;
      END
   END n_132892

   PIN n_132893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.066 0.163 118.094 ;
      END
   END n_132893

   PIN n_132961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.874 122.077 45.902 122.24 ;
      END
   END n_132961

   PIN n_132962
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.81 122.077 45.838 122.24 ;
      END
   END n_132962

   PIN n_133201
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 114.61 0.163 114.638 ;
      END
   END n_133201

   PIN n_133273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 83.314 0.163 83.342 ;
      END
   END n_133273

   PIN n_133287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 83.378 0.163 83.406 ;
      END
   END n_133287

   PIN n_133303
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 111.218 122.077 111.246 122.24 ;
      END
   END n_133303

   PIN n_133427
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.546 122.077 26.574 122.24 ;
      END
   END n_133427

   PIN n_133450
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.378 122.077 307.406 122.24 ;
      END
   END n_133450

   PIN n_133506
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 56.37 0.163 56.398 ;
      END
   END n_133506

   PIN n_133858
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 287.73 122.077 287.758 122.24 ;
      END
   END n_133858

   PIN n_133861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.618 0.163 101.646 ;
      END
   END n_133861

   PIN n_133939
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.314 122.077 307.342 122.24 ;
      END
   END n_133939

   PIN n_134000
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 83.25 0.163 83.278 ;
      END
   END n_134000

   PIN n_134256
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 303.09 122.077 303.118 122.24 ;
      END
   END n_134256

   PIN n_134400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 97.394 0.163 97.422 ;
      END
   END n_134400

   PIN n_134706
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 283.89 122.077 283.918 122.24 ;
      END
   END n_134706

   PIN n_134708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.458 122.077 169.486 122.24 ;
      END
   END n_134708

   PIN n_134825
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.194 0.163 86.222 ;
      END
   END n_134825

   PIN n_134924
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.426 0.163 101.454 ;
      END
   END n_134924

   PIN n_134992
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 7.73 122.077 7.758 122.24 ;
      END
   END n_134992

   PIN n_135296
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 280.114 122.077 280.142 122.24 ;
      END
   END n_135296

   PIN n_135308
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.13 0.163 86.158 ;
      END
   END n_135308

   PIN n_135370
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.306 122.077 176.334 122.24 ;
      END
   END n_135370

   PIN n_135438
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.17 0.163 109.198 ;
      END
   END n_135438

   PIN n_135524
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.034 0.163 90.062 ;
      END
   END n_135524

   PIN n_135528
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.322 122.077 54.35 122.24 ;
      END
   END n_135528

   PIN n_135704
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.154 122.077 311.182 122.24 ;
      END
   END n_135704

   PIN n_135859
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.978 0.163 45.006 ;
      END
   END n_135859

   PIN n_135947
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 53.554 122.077 53.582 122.24 ;
      END
   END n_135947

   PIN n_135957
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.146 122.077 60.174 122.24 ;
      END
   END n_135957

   PIN n_136054
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 307.058 122.077 307.086 122.24 ;
      END
   END n_136054

   PIN n_136077
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 295.41 122.077 295.438 122.24 ;
      END
   END n_136077

   PIN n_136078
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 253.234 122.077 253.262 122.24 ;
      END
   END n_136078

   PIN n_136095
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.786 122.077 172.814 122.24 ;
      END
   END n_136095

   PIN n_136295
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 283.954 122.077 283.982 122.24 ;
      END
   END n_136295

   PIN n_136526
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.394 122.077 57.422 122.24 ;
      END
   END n_136526

   PIN n_136551
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 280.114 122.077 280.142 122.24 ;
      END
   END n_136551

   PIN n_136552
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 280.05 122.077 280.078 122.24 ;
      END
   END n_136552

   PIN n_136555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 276.274 122.077 276.302 122.24 ;
      END
   END n_136555

   PIN n_136727
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 273.778 122.077 273.806 122.24 ;
      END
   END n_136727

   PIN n_136754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 279.986 122.077 280.014 122.24 ;
      END
   END n_136754

   PIN n_136800
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 306.994 122.077 307.022 122.24 ;
      END
   END n_136800

   PIN n_136807
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 291.634 122.077 291.662 122.24 ;
      END
   END n_136807

   PIN n_136808
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 291.57 122.077 291.598 122.24 ;
      END
   END n_136808

   PIN n_136922
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.066 122.077 182.094 122.24 ;
      END
   END n_136922

   PIN n_136951
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 283.762 122.077 283.79 122.24 ;
      END
   END n_136951

   PIN n_137637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 57.394 122.077 57.422 122.24 ;
      END
   END n_137637

   PIN n_137650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 276.21 122.077 276.238 122.24 ;
      END
   END n_137650

   PIN n_14254
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.226 122.077 34.254 122.24 ;
      END
   END n_14254

   PIN n_14255
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.482 122.077 26.51 122.24 ;
      END
   END n_14255

   PIN n_14287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.058 0.163 67.086 ;
      END
   END n_14287

   PIN n_142906
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 110.194 0.163 110.222 ;
      END
   END n_142906

   PIN n_142909
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 117.426 0.163 117.454 ;
      END
   END n_142909

   PIN n_143255
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 228.594 122.077 228.622 122.24 ;
      END
   END n_143255

   PIN n_143341
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.458 122.077 145.486 122.24 ;
      END
   END n_143341

   PIN n_143721
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.362 0.163 101.39 ;
      END
   END n_143721

   PIN n_143848
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 70.962 0.163 70.99 ;
      END
   END n_143848

   PIN n_144235
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 102.066 0.163 102.094 ;
      END
   END n_144235

   PIN n_144239
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 20.658 0.163 20.686 ;
      END
   END n_144239

   PIN n_144318
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 67.25 0.163 67.278 ;
      END
   END n_144318

   PIN n_14452
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 260.85 122.077 260.878 122.24 ;
      END
   END n_14452

   PIN n_14557
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.338 0.163 12.366 ;
      END
   END n_14557

   PIN n_14659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 214.642 122.077 214.67 122.24 ;
      END
   END n_14659

   PIN n_14956
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 219.506 122.077 219.534 122.24 ;
      END
   END n_14956

   PIN n_15206
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 105.65 0.163 105.678 ;
      END
   END n_15206

   PIN n_15462
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 219.378 122.077 219.406 122.24 ;
      END
   END n_15462

   PIN n_16034
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 242.354 122.077 242.382 122.24 ;
      END
   END n_16034

   PIN n_16166
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.234 0.163 109.262 ;
      END
   END n_16166

   PIN n_16255
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.434 122.077 176.462 122.24 ;
      END
   END n_16255

   PIN n_16364
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 7.794 122.077 7.822 122.24 ;
      END
   END n_16364

   PIN n_16366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 283.89 122.077 283.918 122.24 ;
      END
   END n_16366

   PIN n_16486
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 93.682 0.163 93.71 ;
      END
   END n_16486

   PIN n_17494
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 77.682 0.163 77.71 ;
      END
   END n_17494

   PIN n_17661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.354 0.163 114.382 ;
      END
   END n_17661

   PIN n_17796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.29 0.163 114.318 ;
      END
   END n_17796

   PIN n_18022
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 237.938 122.077 237.966 122.24 ;
      END
   END n_18022

   PIN n_18128
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 177.714 122.077 177.742 122.24 ;
      END
   END n_18128

   PIN n_18199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.562 122.077 224.59 122.24 ;
      END
   END n_18199

   PIN n_18869
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.778 122.077 145.806 122.24 ;
      END
   END n_18869

   PIN n_18877
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 283.826 122.077 283.854 122.24 ;
      END
   END n_18877

   PIN n_18948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.37 122.077 176.398 122.24 ;
      END
   END n_18948

   PIN n_18989
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.97 122.077 145.998 122.24 ;
      END
   END n_18989

   PIN n_19350
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.458 122.077 241.486 122.24 ;
      END
   END n_19350

   PIN n_19373
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 183.666 122.077 183.694 122.24 ;
      END
   END n_19373

   PIN n_19607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 134.194 122.077 134.222 122.24 ;
      END
   END n_19607

   PIN n_19629
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 172.594 122.077 172.622 122.24 ;
      END
   END n_19629

   PIN n_19657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 172.53 122.077 172.558 122.24 ;
      END
   END n_19657

   PIN n_19681
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 141.746 122.077 141.774 122.24 ;
      END
   END n_19681

   PIN n_19914
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.514 122.077 126.542 122.24 ;
      END
   END n_19914

   PIN n_19971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 172.53 122.077 172.558 122.24 ;
      END
   END n_19971

   PIN n_19983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 98.034 0.163 98.062 ;
      END
   END n_19983

   PIN n_20006
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 130.418 122.077 130.446 122.24 ;
      END
   END n_20006

   PIN n_20085
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 187.89 122.077 187.918 122.24 ;
      END
   END n_20085

   PIN n_20090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 189.618 122.077 189.646 122.24 ;
      END
   END n_20090

   PIN n_20275
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 283.826 122.077 283.854 122.24 ;
      END
   END n_20275

   PIN n_20413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.986 122.077 88.014 122.24 ;
      END
   END n_20413

   PIN n_20639
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 97.714 0.163 97.742 ;
      END
   END n_20639

   PIN n_20872
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.234 122.077 157.262 122.24 ;
      END
   END n_20872

   PIN n_21109
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 97.97 0.163 97.998 ;
      END
   END n_21109

   PIN n_21129
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 241.202 122.077 241.23 122.24 ;
      END
   END n_21129

   PIN n_21187
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.778 0.163 113.806 ;
      END
   END n_21187

   PIN n_21414
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 198.77 122.077 198.798 122.24 ;
      END
   END n_21414

   PIN n_21637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 114.93 122.077 114.958 122.24 ;
      END
   END n_21637

   PIN n_21657
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 149.49 122.077 149.518 122.24 ;
      END
   END n_21657

   PIN n_21680
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 196.914 122.077 196.942 122.24 ;
      END
   END n_21680

   PIN n_21703
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 114.098 0.163 114.126 ;
      END
   END n_21703

   PIN n_21708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 98.418 0.163 98.446 ;
      END
   END n_21708

   PIN n_21709
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 145.906 122.077 145.934 122.24 ;
      END
   END n_21709

   PIN n_21771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.594 122.077 76.622 122.24 ;
      END
   END n_21771

   PIN n_21806
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.218 122.077 79.246 122.24 ;
      END
   END n_21806

   PIN n_22159
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.594 122.077 76.622 122.24 ;
      END
   END n_22159

   PIN n_22224
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 109.426 0.163 109.454 ;
      END
   END n_22224

   PIN n_22231
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 93.618 0.163 93.646 ;
      END
   END n_22231

   PIN n_22243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 91.506 122.077 91.534 122.24 ;
      END
   END n_22243

   PIN n_22795
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.586 0.163 105.614 ;
      END
   END n_22795

   PIN n_22822
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 145.714 122.077 145.742 122.24 ;
      END
   END n_22822

   PIN n_23394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 214.258 122.077 214.286 122.24 ;
      END
   END n_23394

   PIN n_23404
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 141.938 122.077 141.966 122.24 ;
      END
   END n_23404

   PIN n_23460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 195.506 122.077 195.534 122.24 ;
      END
   END n_23460

   PIN n_24014
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.546 122.077 122.574 122.24 ;
      END
   END n_24014

   PIN n_24074
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 229.426 122.077 229.454 122.24 ;
      END
   END n_24074

   PIN n_24124
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 224.69 122.077 224.718 122.24 ;
      END
   END n_24124

   PIN n_24141
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.482 122.077 218.51 122.24 ;
      END
   END n_24141

   PIN n_24645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 126.514 122.077 126.542 122.24 ;
      END
   END n_24645

   PIN n_24723
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 111.09 122.077 111.118 122.24 ;
      END
   END n_24723

   PIN n_24774
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 248.498 122.077 248.526 122.24 ;
      END
   END n_24774

   PIN n_25460
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 113.394 0.163 113.422 ;
      END
   END n_25460

   PIN n_26642
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 207.602 122.077 207.63 122.24 ;
      END
   END n_26642

   PIN n_28886
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 295.474 122.077 295.502 122.24 ;
      END
   END n_28886

   PIN n_31620
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.898 122.077 22.926 122.24 ;
      END
   END n_31620

   PIN n_31789
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 113.394 313.394 113.422 ;
      END
   END n_31789

   PIN n_32482
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 82.61 313.394 82.638 ;
      END
   END n_32482

   PIN n_32483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 313.23 105.65 313.394 105.678 ;
      END
   END n_32483

   PIN n_32637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.298 0.163 117.326 ;
      END
   END n_32637

   PIN n_32919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.154 122.077 15.182 122.24 ;
      END
   END n_32919

   PIN n_32920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.026 122.077 15.054 122.24 ;
      END
   END n_32920

   PIN n_32934
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.002 0.163 86.03 ;
      END
   END n_32934

   PIN n_33003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 86.066 0.163 86.094 ;
      END
   END n_33003

   PIN n_33076
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.69 122.077 72.718 122.24 ;
      END
   END n_33076

   PIN n_33077
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.01 122.077 129.038 122.24 ;
      END
   END n_33077

   PIN n_33264
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 287.666 122.077 287.694 122.24 ;
      END
   END n_33264

   PIN n_33268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.09 122.077 311.118 122.24 ;
      END
   END n_33268

   PIN n_33473
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 82.93 0.163 82.958 ;
      END
   END n_33473

   PIN n_33483
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.938 0.163 101.966 ;
      END
   END n_33483

   PIN n_33921
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.554 0.163 101.582 ;
      END
   END n_33921

   PIN n_33953
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.97 122.077 41.998 122.24 ;
      END
   END n_33953

   PIN n_34366
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.098 122.077 42.126 122.24 ;
      END
   END n_34366

   PIN n_34708
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 117.106 0.163 117.134 ;
      END
   END n_34708

   PIN n_34720
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.018 122.077 124.046 122.24 ;
      END
   END n_34720

   PIN n_35010
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.146 122.077 20.174 122.24 ;
      END
   END n_35010

   PIN n_35016
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.234 122.077 61.262 122.24 ;
      END
   END n_35016

   PIN n_35029
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.202 122.077 33.23 122.24 ;
      END
   END n_35029

   PIN n_35032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.034 122.077 34.062 122.24 ;
      END
   END n_35032

   PIN n_35033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.354 122.077 34.382 122.24 ;
      END
   END n_35033

   PIN n_35070
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 291.506 122.077 291.534 122.24 ;
      END
   END n_35070

   PIN n_35739
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.938 122.077 45.966 122.24 ;
      END
   END n_35739

   PIN n_36449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.33 0.163 17.358 ;
      END
   END n_36449

   PIN n_3711
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 101.49 0.163 101.518 ;
      END
   END n_3711

   PIN n_3868
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 86.194 0.163 86.222 ;
      END
   END n_3868

   PIN n_39087
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.554 0.163 117.582 ;
      END
   END n_39087

   PIN n_39278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 94.514 0.163 94.542 ;
      END
   END n_39278

   PIN n_3945
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 311.026 122.077 311.054 122.24 ;
      END
   END n_3945

   PIN n_39484
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 118.002 0.163 118.03 ;
      END
   END n_39484

   PIN n_39485
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 117.938 0.163 117.966 ;
      END
   END n_39485

   PIN n_41711
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 272.498 122.077 272.526 122.24 ;
      END
   END n_41711

   PIN n_4199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.042 122.077 61.07 122.24 ;
      END
   END n_4199

   PIN n_5193
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.306 122.077 80.334 122.24 ;
      END
   END n_5193

   PIN n_5196
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.682 0.163 101.71 ;
      END
   END n_5196

   PIN n_5565
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.946 122.077 64.974 122.24 ;
      END
   END n_5565

   PIN n_6522
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.738 0.163 90.766 ;
      END
   END n_6522

   PIN n_6525
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 105.97 0.163 105.998 ;
      END
   END n_6525

   PIN n_6542
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 108.914 0.163 108.942 ;
      END
   END n_6542

   PIN n_6619
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 110.962 122.077 110.99 122.24 ;
      END
   END n_6619

   PIN n_6693
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.362 0.163 53.39 ;
      END
   END n_6693

   PIN n_6697
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 78.45 0.163 78.478 ;
      END
   END n_6697

   PIN n_6937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 63.474 0.163 63.502 ;
      END
   END n_6937

   PIN n_7273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 176.306 122.077 176.334 122.24 ;
      END
   END n_7273

   PIN n_8119
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 101.49 0.163 101.518 ;
      END
   END n_8119

   PIN n_8247
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.258 0.163 62.286 ;
      END
   END n_8247

   PIN n_8343
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 67.378 0.163 67.406 ;
      END
   END n_8343

   PIN n_8387
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 130.226 122.077 130.254 122.24 ;
      END
   END n_8387

   PIN n_890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 90.418 0.163 90.446 ;
      END
   END n_890

   PIN n_912
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 40.37 0.163 40.398 ;
      END
   END n_912

   PIN n_9132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 219.57 122.077 219.598 122.24 ;
      END
   END n_9132

   PIN n_9798
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.666 0.163 55.694 ;
      END
   END n_9798

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 313.394 122.24 ;
      LAYER V1 ;
         RECT 0.0 0.0 313.394 122.24 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 313.394 122.24 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 313.394 122.24 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 313.394 122.24 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 313.394 122.24 ;
      LAYER M1 ;
         RECT 0.0 0.0 313.394 122.24 ;
   END
END h0_mgc_matrix_mult_b

MACRO h5_mgc_fft_a
   CLASS BLOCK ;
   FOREIGN h5 ;
   ORIGIN 0 0 ;
   SIZE 97.024 BY 46.08 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1102_rst
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.866 0.0 90.894 0.163 ;
      END
   END FE_OFN1102_rst

   PIN FE_OFN267_n_4280
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.474 45.998 79.502 46.08 ;
      END
   END FE_OFN267_n_4280

   PIN FE_OFN827_n_3772
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 44.722 97.024 44.75 ;
      END
   END FE_OFN827_n_3772

   PIN FE_OFN829_n_8424
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.114 45.917 88.142 46.08 ;
      END
   END FE_OFN829_n_8424

   PIN n_10129
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.578 0.163 38.606 ;
      END
   END n_10129

   PIN n_10572
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.442 0.163 43.47 ;
      END
   END n_10572

   PIN n_10650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.17 0.0 37.198 0.163 ;
      END
   END n_10650

   PIN n_10952
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.874 0.0 29.902 0.163 ;
      END
   END n_10952

   PIN n_10953
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.634 0.0 27.662 0.163 ;
      END
   END n_10953

   PIN n_12076
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.21 45.917 28.238 46.08 ;
      END
   END n_12076

   PIN n_12100
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.666 0.0 31.694 0.163 ;
      END
   END n_12100

   PIN n_12221
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.802 0.0 34.83 0.163 ;
      END
   END n_12221

   PIN n_1247
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 78.962 45.917 78.99 46.08 ;
      END
   END n_1247

   PIN n_12608
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.442 0.163 27.47 ;
      END
   END n_12608

   PIN n_12826
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.49 45.917 29.518 46.08 ;
      END
   END n_12826

   PIN n_13290
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.93 0.0 10.958 0.163 ;
      END
   END n_13290

   PIN n_13898
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.25 0.163 27.278 ;
      END
   END n_13898

   PIN n_14243
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.57 0.0 27.598 0.163 ;
      END
   END n_14243

   PIN n_14244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.554 0.0 29.582 0.163 ;
      END
   END n_14244

   PIN n_14522
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.202 45.917 81.23 46.08 ;
      END
   END n_14522

   PIN n_14855
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.394 0.0 33.422 0.163 ;
      END
   END n_14855

   PIN n_14856
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.33 0.0 33.358 0.163 ;
      END
   END n_14856

   PIN n_1487
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 22.834 97.024 22.862 ;
      END
   END n_1487

   PIN n_15005
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 38.386 97.024 38.414 ;
      END
   END n_15005

   PIN n_15031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.818 0.0 24.846 0.163 ;
      END
   END n_15031

   PIN n_15092
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.506 0.0 27.534 0.163 ;
      END
   END n_15092

   PIN n_15377
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.45 0.0 30.478 0.163 ;
      END
   END n_15377

   PIN n_1591
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.298 45.917 85.326 46.08 ;
      END
   END n_1591

   PIN n_15967
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 35.954 97.024 35.982 ;
      END
   END n_15967

   PIN n_16054
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.97 0.0 25.998 0.163 ;
      END
   END n_16054

   PIN n_16555
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.706 0.163 22.734 ;
      END
   END n_16555

   PIN n_16749
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.77 0.163 22.798 ;
      END
   END n_16749

   PIN n_16770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.034 0.0 26.062 0.163 ;
      END
   END n_16770

   PIN n_17130
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.138 0.0 17.166 0.163 ;
      END
   END n_17130

   PIN n_17673
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.146 0.0 28.174 0.163 ;
      END
   END n_17673

   PIN n_19031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.306 0.163 24.334 ;
      END
   END n_19031

   PIN n_19333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.77 0.0 14.798 0.163 ;
      END
   END n_19333

   PIN n_19372
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.898 0.163 22.926 ;
      END
   END n_19372

   PIN n_20390
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 4.274 97.024 4.302 ;
      END
   END n_20390

   PIN n_2339
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.538 45.917 15.566 46.08 ;
      END
   END n_2339

   PIN n_23513
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 12.85 97.024 12.878 ;
      END
   END n_23513

   PIN n_24465
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.178 0.0 72.206 0.163 ;
      END
   END n_24465

   PIN n_25465
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.01 45.917 73.038 46.08 ;
      END
   END n_25465

   PIN n_26031
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.258 45.917 70.286 46.08 ;
      END
   END n_26031

   PIN n_27335
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 2.674 97.024 2.702 ;
      END
   END n_27335

   PIN n_28336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 12.786 97.024 12.814 ;
      END
   END n_28336

   PIN n_28551
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.562 45.917 48.59 46.08 ;
      END
   END n_28551

   PIN n_28552
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.498 45.917 48.526 46.08 ;
      END
   END n_28552

   PIN n_28705
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 2.61 97.024 2.638 ;
      END
   END n_28705

   PIN n_29060
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 4.338 97.024 4.366 ;
      END
   END n_29060

   PIN n_29114
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.17 45.917 85.198 46.08 ;
      END
   END n_29114

   PIN n_29356
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 38.322 97.024 38.35 ;
      END
   END n_29356

   PIN n_29588
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.394 45.917 73.422 46.08 ;
      END
   END n_29588

   PIN n_29605
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.658 45.917 76.686 46.08 ;
      END
   END n_29605

   PIN n_2970
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.81 45.917 21.838 46.08 ;
      END
   END n_2970

   PIN n_3176
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 43.442 97.024 43.47 ;
      END
   END n_3176

   PIN n_3798
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.874 45.917 21.902 46.08 ;
      END
   END n_3798

   PIN n_3802
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 21.938 45.917 21.966 46.08 ;
      END
   END n_3802

   PIN n_3839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.05 45.917 16.078 46.08 ;
      END
   END n_3839

   PIN n_4058
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.93 45.917 18.958 46.08 ;
      END
   END n_4058

   PIN n_4072
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.778 45.917 25.806 46.08 ;
      END
   END n_4072

   PIN n_5262
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.234 45.917 85.262 46.08 ;
      END
   END n_5262

   PIN n_5327
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.106 45.917 85.134 46.08 ;
      END
   END n_5327

   PIN n_5340
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.562 45.917 16.59 46.08 ;
      END
   END n_5340

   PIN n_5341
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.234 45.917 13.262 46.08 ;
      END
   END n_5341

   PIN n_5519
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.41 45.917 79.438 46.08 ;
      END
   END n_5519

   PIN n_6244
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.258 0.163 30.286 ;
      END
   END n_6244

   PIN n_6256
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.882 45.917 24.91 46.08 ;
      END
   END n_6256

   PIN n_6595
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.074 0.0 33.102 0.163 ;
      END
   END n_6595

   PIN n_6979
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.13 0.163 30.158 ;
      END
   END n_6979

   PIN n_6987
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.194 0.163 30.222 ;
      END
   END n_6987

   PIN n_7017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.714 45.917 1.742 46.08 ;
      END
   END n_7017

   PIN n_7224
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.154 45.917 39.182 46.08 ;
      END
   END n_7224

   PIN n_7237
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 30.194 97.024 30.222 ;
      END
   END n_7237

   PIN n_7274
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.57 45.917 19.598 46.08 ;
      END
   END n_7274

   PIN n_7311
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.594 45.917 76.622 46.08 ;
      END
   END n_7311

   PIN n_8443
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.586 45.917 25.614 46.08 ;
      END
   END n_8443

   PIN n_8444
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.754 45.917 24.782 46.08 ;
      END
   END n_8444

   PIN n_9230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.29 0.163 34.318 ;
      END
   END n_9230

   PIN n_9350
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.386 0.163 38.414 ;
      END
   END n_9350

   PIN n_9351
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.45 0.163 38.478 ;
      END
   END n_9351

   PIN n_9728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.314 0.163 27.342 ;
      END
   END n_9728

   PIN n_9943
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.106 45.917 37.134 46.08 ;
      END
   END n_9943

   PIN x_out_21_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 24.37 97.024 24.398 ;
      END
   END x_out_21_1

   PIN x_out_21_22
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 35.89 97.024 35.918 ;
      END
   END x_out_21_22

   PIN x_out_21_23
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 21.49 97.024 21.518 ;
      END
   END x_out_21_23

   PIN x_out_21_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 38.834 97.024 38.862 ;
      END
   END x_out_21_24

   PIN x_out_21_25
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 30.002 97.024 30.03 ;
      END
   END x_out_21_25

   PIN x_out_21_26
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 19.826 97.024 19.854 ;
      END
   END x_out_21_26

   PIN x_out_25_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 12.914 97.024 12.942 ;
      END
   END x_out_25_29

   PIN x_out_25_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 7.09 97.024 7.118 ;
      END
   END x_out_25_30

   PIN x_out_53_22
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 27.122 97.024 27.15 ;
      END
   END x_out_53_22

   PIN x_out_53_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 35.89 97.024 35.918 ;
      END
   END x_out_53_24

   PIN x_out_53_25
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 30.13 97.024 30.158 ;
      END
   END x_out_53_25

   PIN x_out_53_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 35.826 97.024 35.854 ;
      END
   END x_out_53_28

   PIN x_out_55_14
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 38.77 97.024 38.798 ;
      END
   END x_out_55_14

   PIN x_out_57_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 29.874 97.024 29.902 ;
      END
   END x_out_57_29

   PIN x_out_57_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 27.058 97.024 27.086 ;
      END
   END x_out_57_30

   PIN x_out_5_13
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 33.266 97.024 33.294 ;
      END
   END x_out_5_13

   PIN FE_OFN1171_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 93.362 0.0 93.39 0.163 ;
      END
   END FE_OFN1171_n_4860

   PIN FE_OFN1264_n_29354
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.994 45.917 91.022 46.08 ;
      END
   END FE_OFN1264_n_29354

   PIN FE_OFN184_n_29402
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 33.202 97.024 33.23 ;
      END
   END FE_OFN184_n_29402

   PIN FE_OFN248_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.942 26.93 97.024 26.958 ;
      END
   END FE_OFN248_n_4162

   PIN FE_OFN261_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.77 45.917 30.798 46.08 ;
      END
   END FE_OFN261_n_4280

   PIN FE_OFN300_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 81.394 45.998 81.422 46.08 ;
      END
   END FE_OFN300_n_3069

   PIN FE_OFN303_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.746 0.0 77.774 0.082 ;
      END
   END FE_OFN303_n_3069

   PIN FE_OFN308_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.426 45.917 85.454 46.08 ;
      END
   END FE_OFN308_n_3069

   PIN FE_OFN326_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.594 45.998 76.622 46.08 ;
      END
   END FE_OFN326_n_4860

   PIN FE_OFN347_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.942 22.45 97.024 22.478 ;
      END
   END FE_OFN347_n_4860

   PIN FE_OFN35_n_15183
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 61.618 45.917 61.646 46.08 ;
      END
   END FE_OFN35_n_15183

   PIN FE_OFN400_n_28303
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 84.978 0.0 85.006 0.082 ;
      END
   END FE_OFN400_n_28303

   PIN FE_OFN56_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 33.266 0.082 33.294 ;
      END
   END FE_OFN56_n_27012

   PIN FE_OFN89_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 84.402 45.998 84.43 46.08 ;
      END
   END FE_OFN89_n_27449

   PIN FE_OFN90_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.942 33.522 97.024 33.55 ;
      END
   END FE_OFN90_n_27449

   PIN FE_OFN91_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.658 45.917 84.686 46.08 ;
      END
   END FE_OFN91_n_27449

   PIN FE_OFN92_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 91.058 45.998 91.086 46.08 ;
      END
   END FE_OFN92_n_27449

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.942 38.514 97.024 38.542 ;
      END
   END ispd_clk

   PIN n_10128
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.514 0.163 38.542 ;
      END
   END n_10128

   PIN n_14910
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.378 0.163 27.406 ;
      END
   END n_14910

   PIN n_15268
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 22.642 97.024 22.67 ;
      END
   END n_15268

   PIN n_15269
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 24.306 97.024 24.334 ;
      END
   END n_15269

   PIN n_15378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.282 0.0 23.31 0.163 ;
      END
   END n_15378

   PIN n_15877
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 24.754 0.0 24.782 0.163 ;
      END
   END n_15877

   PIN n_15878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.13 0.0 22.158 0.163 ;
      END
   END n_15878

   PIN n_15922
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 17.842 97.024 17.87 ;
      END
   END n_15922

   PIN n_17184
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 22.77 97.024 22.798 ;
      END
   END n_17184

   PIN n_17474
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.714 0.0 17.742 0.163 ;
      END
   END n_17474

   PIN n_17671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.378 0.0 27.406 0.163 ;
      END
   END n_17671

   PIN n_17672
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.21 0.0 28.238 0.163 ;
      END
   END n_17672

   PIN n_19032
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.242 0.163 24.27 ;
      END
   END n_19032

   PIN n_21830
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.338 0.0 92.366 0.163 ;
      END
   END n_21830

   PIN n_22019
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 93.17 45.998 93.198 46.08 ;
      END
   END n_22019

   PIN n_22492
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 92.274 0.0 92.302 0.163 ;
      END
   END n_22492

   PIN n_23182
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 12.786 0.163 12.814 ;
      END
   END n_23182

   PIN n_2343
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 21.298 97.024 21.326 ;
      END
   END n_2343

   PIN n_237
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 17.906 97.024 17.934 ;
      END
   END n_237

   PIN n_23813
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 9.266 45.998 9.294 46.08 ;
      END
   END n_23813

   PIN n_24424
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.298 45.917 13.326 46.08 ;
      END
   END n_24424

   PIN n_24865
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.002 45.917 22.03 46.08 ;
      END
   END n_24865

   PIN n_26084
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.994 45.917 19.022 46.08 ;
      END
   END n_26084

   PIN n_26271
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.954 0.163 35.982 ;
      END
   END n_26271

   PIN n_26570
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.322 0.163 38.35 ;
      END
   END n_26570

   PIN n_27334
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 2.546 97.024 2.574 ;
      END
   END n_27334

   PIN n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.154 45.998 39.182 46.08 ;
      END
   END n_27449

   PIN n_28550
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.538 45.917 47.566 46.08 ;
      END
   END n_28550

   PIN n_28597
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.034 45.917 90.062 46.08 ;
      END
   END n_28597

   PIN n_29046
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.946 45.998 40.974 46.08 ;
      END
   END n_29046

   PIN n_29068
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.73 45.917 31.758 46.08 ;
      END
   END n_29068

   PIN n_29126
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.266 45.917 25.294 46.08 ;
      END
   END n_29126

   PIN n_29261
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.942 33.394 97.024 33.422 ;
      END
   END n_29261

   PIN n_29664
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 13.17 45.998 13.198 46.08 ;
      END
   END n_29664

   PIN n_29683
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.942 44.594 97.024 44.622 ;
      END
   END n_29683

   PIN n_5003
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.466 45.917 76.494 46.08 ;
      END
   END n_5003

   PIN n_5445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.266 45.917 25.294 46.08 ;
      END
   END n_5445

   PIN n_546
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.01 45.917 41.038 46.08 ;
      END
   END n_546

   PIN n_7214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 19.762 97.024 19.79 ;
      END
   END n_7214

   PIN n_8671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.626 45.917 16.654 46.08 ;
      END
   END n_8671

   PIN rst
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 90.93 45.998 90.958 46.08 ;
      END
   END rst

   PIN x_in_39_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 22.578 97.024 22.606 ;
      END
   END x_in_39_13

   PIN x_in_39_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 21.618 97.024 21.646 ;
      END
   END x_in_39_14

   PIN x_in_39_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 22.706 97.024 22.734 ;
      END
   END x_in_39_15

   PIN x_in_42_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.41 0.0 23.438 0.163 ;
      END
   END x_in_42_1

   PIN x_in_42_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 10.802 97.024 10.83 ;
      END
   END x_in_42_10

   PIN x_in_42_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.594 0.0 76.622 0.163 ;
      END
   END x_in_42_11

   PIN x_in_42_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 24.242 97.024 24.27 ;
      END
   END x_in_42_12

   PIN x_in_42_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 30.514 97.024 30.542 ;
      END
   END x_in_42_13

   PIN x_in_42_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 30.45 97.024 30.478 ;
      END
   END x_in_42_14

   PIN x_in_42_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 33.522 97.024 33.55 ;
      END
   END x_in_42_15

   PIN x_in_43_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 7.666 97.024 7.694 ;
      END
   END x_in_43_0

   PIN x_in_43_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 15.794 97.024 15.822 ;
      END
   END x_in_43_1

   PIN x_in_43_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 30.386 97.024 30.414 ;
      END
   END x_in_43_10

   PIN x_in_43_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.834 45.998 22.862 46.08 ;
      END
   END x_in_43_11

   PIN x_in_43_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 27.314 97.024 27.342 ;
      END
   END x_in_43_12

   PIN x_in_43_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.866 45.917 50.894 46.08 ;
      END
   END x_in_43_13

   PIN x_in_43_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.602 45.917 55.63 46.08 ;
      END
   END x_in_43_14

   PIN x_in_43_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 36.082 97.024 36.11 ;
      END
   END x_in_43_15

   PIN x_in_43_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 7.282 97.024 7.31 ;
      END
   END x_in_43_2

   PIN x_in_43_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 10.93 97.024 10.958 ;
      END
   END x_in_43_3

   PIN x_in_43_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 54.45 45.998 54.478 46.08 ;
      END
   END x_in_43_4

   PIN x_in_43_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.942 24.754 97.024 24.782 ;
      END
   END x_in_43_5

   PIN x_in_43_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 19.89 97.024 19.918 ;
      END
   END x_in_43_6

   PIN x_in_43_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.861 24.626 97.024 24.654 ;
      END
   END x_in_43_7

   PIN x_in_43_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.942 22.066 97.024 22.094 ;
      END
   END x_in_43_8

   PIN x_in_43_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.942 27.378 97.024 27.406 ;
      END
   END x_in_43_9

   PIN x_out_21_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.354 45.917 82.382 46.08 ;
      END
   END x_out_21_15

   PIN x_out_21_20
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 87.09 45.917 87.118 46.08 ;
      END
   END x_out_21_20

   PIN x_out_21_21
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.026 45.917 79.054 46.08 ;
      END
   END x_out_21_21

   PIN x_out_25_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.861 22.898 97.024 22.926 ;
      END
   END x_out_25_15

   PIN x_out_53_26
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.418 45.917 82.446 46.08 ;
      END
   END x_out_53_26

   PIN x_out_57_31
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.834 0.163 22.862 ;
      END
   END x_out_57_31

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 97.024 46.08 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 97.024 46.08 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 97.024 46.08 ;
      LAYER V1 ;
         RECT 0.0 0.0 97.024 46.08 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 97.024 46.08 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 97.024 46.08 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 97.024 46.08 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 97.024 46.08 ;
      LAYER M1 ;
         RECT 0.0 0.0 97.024 46.08 ;
   END
END h5_mgc_fft_a

MACRO h4_mgc_fft_a
   CLASS BLOCK ;
   FOREIGN h4 ;
   ORIGIN 0 0 ;
   SIZE 99.52 BY 67.84 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN276_n_16893
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 0.946 67.677 0.974 67.84 ;
      END
   END FE_OFN276_n_16893

   PIN FE_OFN282_n_7349
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 46.642 0.163 46.67 ;
      END
   END FE_OFN282_n_7349

   PIN FE_OFN339_n_4860
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.594 0.163 60.622 ;
      END
   END FE_OFN339_n_4860

   PIN FE_OFN352_n_4860
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.69 0.082 48.718 ;
      END
   END FE_OFN352_n_4860

   PIN n_10750
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.314 0.163 27.342 ;
      END
   END n_10750

   PIN n_12144
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 55.538 67.677 55.566 67.84 ;
      END
   END n_12144

   PIN n_1289
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 44.658 67.677 44.686 67.84 ;
      END
   END n_1289

   PIN n_13764
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 64.882 0.163 64.91 ;
      END
   END n_13764

   PIN n_14521
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.154 67.677 63.182 67.84 ;
      END
   END n_14521

   PIN n_14885
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 59.186 0.163 59.214 ;
      END
   END n_14885

   PIN n_15325
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.794 0.163 39.822 ;
      END
   END n_15325

   PIN n_15907
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.122 0.163 59.15 ;
      END
   END n_15907

   PIN n_16753
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.53 0.163 44.558 ;
      END
   END n_16753

   PIN n_16798
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.482 0.163 50.51 ;
      END
   END n_16798

   PIN n_17335
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.066 0.163 62.094 ;
      END
   END n_17335

   PIN n_17762
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.074 0.163 65.102 ;
      END
   END n_17762

   PIN n_17906
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.658 0.163 60.686 ;
      END
   END n_17906

   PIN n_17993
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.322 0.163 62.35 ;
      END
   END n_17993

   PIN n_18103
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.17 0.163 37.198 ;
      END
   END n_18103

   PIN n_18127
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.034 0.163 42.062 ;
      END
   END n_18127

   PIN n_18128
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.97 0.163 41.998 ;
      END
   END n_18128

   PIN n_18481
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.946 0.163 64.974 ;
      END
   END n_18481

   PIN n_18575
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.234 0.163 37.262 ;
      END
   END n_18575

   PIN n_1865
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.41 67.677 39.438 67.84 ;
      END
   END n_1865

   PIN n_18833
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.098 0.163 42.126 ;
      END
   END n_18833

   PIN n_18835
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.906 0.163 41.934 ;
      END
   END n_18835

   PIN n_19121
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.594 0.163 60.622 ;
      END
   END n_19121

   PIN n_19140
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.882 0.163 64.91 ;
      END
   END n_19140

   PIN n_19235
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 62.258 0.163 62.286 ;
      END
   END n_19235

   PIN n_19322
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.826 0.163 27.854 ;
      END
   END n_19322

   PIN n_19382
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.61 0.163 18.638 ;
      END
   END n_19382

   PIN n_19891
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.594 0.163 44.622 ;
      END
   END n_19891

   PIN n_19966
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.01 0.163 65.038 ;
      END
   END n_19966

   PIN n_20233
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.722 0.163 44.75 ;
      END
   END n_20233

   PIN n_20283
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.186 0.163 59.214 ;
      END
   END n_20283

   PIN n_20288
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.698 0.163 51.726 ;
      END
   END n_20288

   PIN n_20344
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.642 0.163 30.67 ;
      END
   END n_20344

   PIN n_20690
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 64.946 0.163 64.974 ;
      END
   END n_20690

   PIN n_20766
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.05 0.163 56.078 ;
      END
   END n_20766

   PIN n_21207
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.818 0.163 64.846 ;
      END
   END n_21207

   PIN n_21332
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.378 0.163 27.406 ;
      END
   END n_21332

   PIN n_21382
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.514 67.677 14.542 67.84 ;
      END
   END n_21382

   PIN n_21383
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.794 67.677 15.822 67.84 ;
      END
   END n_21383

   PIN n_21442
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 56.242 0.163 56.27 ;
      END
   END n_21442

   PIN n_21523
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.362 0.163 37.39 ;
      END
   END n_21523

   PIN n_22114
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.49 0.163 53.518 ;
      END
   END n_22114

   PIN n_22537
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.106 0.163 37.134 ;
      END
   END n_22537

   PIN n_22682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.386 0.163 62.414 ;
      END
   END n_22682

   PIN n_22691
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.53 0.163 60.558 ;
      END
   END n_22691

   PIN n_22799
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.554 0.163 53.582 ;
      END
   END n_22799

   PIN n_23517
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.618 0.163 53.646 ;
      END
   END n_23517

   PIN n_23682
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.138 0.163 65.166 ;
      END
   END n_23682

   PIN n_23683
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.194 0.163 62.222 ;
      END
   END n_23683

   PIN n_23747
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.098 67.677 82.126 67.84 ;
      END
   END n_23747

   PIN n_23770
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.634 0.163 51.662 ;
      END
   END n_23770

   PIN n_23771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.57 0.163 51.598 ;
      END
   END n_23771

   PIN n_24387
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.314 0.163 51.342 ;
      END
   END n_24387

   PIN n_24576
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.746 0.163 53.774 ;
      END
   END n_24576

   PIN n_25009
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.986 0.163 56.014 ;
      END
   END n_25009

   PIN n_25062
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.834 0.163 46.862 ;
      END
   END n_25062

   PIN n_25138
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.434 0.163 32.462 ;
      END
   END n_25138

   PIN n_2520
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.194 0.163 46.222 ;
      END
   END n_2520

   PIN n_2536
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.162 67.677 58.19 67.84 ;
      END
   END n_2536

   PIN n_25410
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.25 0.163 51.278 ;
      END
   END n_25410

   PIN n_25427
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.13 67.677 30.158 67.84 ;
      END
   END n_25427

   PIN n_26633
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 36.21 0.163 36.238 ;
      END
   END n_26633

   PIN n_27097
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.466 67.677 36.494 67.84 ;
      END
   END n_27097

   PIN n_27589
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 36.466 67.677 36.494 67.84 ;
      END
   END n_27589

   PIN n_27724
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.298 0.163 37.326 ;
      END
   END n_27724

   PIN n_27869
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 92.978 67.677 93.006 67.84 ;
      END
   END n_27869

   PIN n_28230
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.418 0.163 50.446 ;
      END
   END n_28230

   PIN n_28326
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.562 67.677 48.59 67.84 ;
      END
   END n_28326

   PIN n_28704
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 51.25 99.52 51.278 ;
      END
   END n_28704

   PIN n_28807
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.282 67.677 31.31 67.84 ;
      END
   END n_28807

   PIN n_28821
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.77 0.163 46.798 ;
      END
   END n_28821

   PIN n_29052
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.354 0.163 10.382 ;
      END
   END n_29052

   PIN n_29059
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 21.81 0.163 21.838 ;
      END
   END n_29059

   PIN n_29152
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.554 0.163 13.582 ;
      END
   END n_29152

   PIN n_29153
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.49 0.163 13.518 ;
      END
   END n_29153

   PIN n_29372
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.418 0.163 10.446 ;
      END
   END n_29372

   PIN n_2947
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.09 0.163 23.118 ;
      END
   END n_2947

   PIN n_2951
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.042 0.163 45.07 ;
      END
   END n_2951

   PIN n_4021
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.258 0.163 46.286 ;
      END
   END n_4021

   PIN n_4881
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.338 0.163 60.366 ;
      END
   END n_4881

   PIN n_5362
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 23.026 0.163 23.054 ;
      END
   END n_5362

   PIN n_5669
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.658 0.163 44.686 ;
      END
   END n_5669

   PIN n_7328
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.106 67.677 45.134 67.84 ;
      END
   END n_7328

   PIN n_8581
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 36.274 0.163 36.302 ;
      END
   END n_8581

   PIN n_9651
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.682 0.163 21.71 ;
      END
   END n_9651

   PIN x_out_22_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 41.842 0.163 41.87 ;
      END
   END x_out_22_12

   PIN x_out_22_13
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 27.57 0.163 27.598 ;
      END
   END x_out_22_13

   PIN x_out_22_14
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 13.106 0.163 13.134 ;
      END
   END x_out_22_14

   PIN x_out_22_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.29 0.163 10.318 ;
      END
   END x_out_22_15

   PIN x_out_22_23
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 50.738 0.163 50.766 ;
      END
   END x_out_22_23

   PIN x_out_22_25
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 53.426 0.163 53.454 ;
      END
   END x_out_22_25

   PIN x_out_22_26
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 53.362 0.163 53.39 ;
      END
   END x_out_22_26

   PIN x_out_22_27
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 60.082 67.677 60.11 67.84 ;
      END
   END x_out_22_27

   PIN x_out_22_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.426 0.163 53.454 ;
      END
   END x_out_22_28

   PIN x_out_27_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 50.674 0.163 50.702 ;
      END
   END x_out_27_0

   PIN x_out_2_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 50.674 0.163 50.702 ;
      END
   END x_out_2_12

   PIN x_out_2_13
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.29 0.163 10.318 ;
      END
   END x_out_2_13

   PIN x_out_2_27
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 59.25 0.163 59.278 ;
      END
   END x_out_2_27

   PIN x_out_2_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 57.65 0.163 57.678 ;
      END
   END x_out_2_28

   PIN x_out_2_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 65.01 0.163 65.038 ;
      END
   END x_out_2_29

   PIN x_out_2_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.018 67.677 28.046 67.84 ;
      END
   END x_out_2_30

   PIN x_out_34_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 41.97 0.163 41.998 ;
      END
   END x_out_34_15

   PIN x_out_34_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 50.866 0.163 50.894 ;
      END
   END x_out_34_28

   PIN x_out_34_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 65.074 0.163 65.102 ;
      END
   END x_out_34_29

   PIN x_out_34_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.394 67.677 33.422 67.84 ;
      END
   END x_out_34_30

   PIN x_out_34_31
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 53.554 0.163 53.582 ;
      END
   END x_out_34_31

   PIN x_out_54_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 51.186 99.52 51.214 ;
      END
   END x_out_54_10

   PIN x_out_54_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 50.61 0.163 50.638 ;
      END
   END x_out_54_11

   PIN x_out_54_14
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 39.858 0.163 39.886 ;
      END
   END x_out_54_14

   PIN x_out_54_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.666 0.163 39.694 ;
      END
   END x_out_54_15

   PIN x_out_54_22
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 24.754 0.163 24.782 ;
      END
   END x_out_54_22

   PIN x_out_54_23
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.986 67.677 48.014 67.84 ;
      END
   END x_out_54_23

   PIN x_out_54_25
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 62.066 0.163 62.094 ;
      END
   END x_out_54_25

   PIN x_out_54_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.402 0.163 60.43 ;
      END
   END x_out_54_29

   PIN x_out_54_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 44.658 0.163 44.686 ;
      END
   END x_out_54_30

   PIN x_out_54_9
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 59.314 99.52 59.342 ;
      END
   END x_out_54_9

   PIN x_out_59_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 53.234 0.163 53.262 ;
      END
   END x_out_59_0

   PIN FE_OFN101_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.858 67.758 47.886 67.84 ;
      END
   END FE_OFN101_n_27449

   PIN FE_OFN105_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 52.722 67.758 52.75 67.84 ;
      END
   END FE_OFN105_n_27449

   PIN FE_OFN1109_rst
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.178 67.758 40.206 67.84 ;
      END
   END FE_OFN1109_rst

   PIN FE_OFN1119_rst
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 47.602 67.758 47.63 67.84 ;
      END
   END FE_OFN1119_rst

   PIN FE_OFN133_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.274 0.082 60.302 ;
      END
   END FE_OFN133_n_27449

   PIN FE_OFN138_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 46.642 0.082 46.67 ;
      END
   END FE_OFN138_n_27449

   PIN FE_OFN175_n_26184
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.058 0.163 59.086 ;
      END
   END FE_OFN175_n_26184

   PIN FE_OFN183_n_29402
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 18.354 99.52 18.382 ;
      END
   END FE_OFN183_n_29402

   PIN FE_OFN212_n_29661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.402 0.163 60.43 ;
      END
   END FE_OFN212_n_29661

   PIN FE_OFN214_n_29687
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.322 67.677 62.35 67.84 ;
      END
   END FE_OFN214_n_29687

   PIN FE_OFN234_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.922 67.758 39.95 67.84 ;
      END
   END FE_OFN234_n_4162

   PIN FE_OFN253_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.914 0.082 44.942 ;
      END
   END FE_OFN253_n_4280

   PIN FE_OFN257_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.438 41.842 99.52 41.87 ;
      END
   END FE_OFN257_n_4280

   PIN FE_OFN271_n_16028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.01 67.677 81.038 67.84 ;
      END
   END FE_OFN271_n_16028

   PIN FE_OFN275_n_16893
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.778 0.163 41.806 ;
      END
   END FE_OFN275_n_16893

   PIN FE_OFN286_n_29266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.586 67.677 33.614 67.84 ;
      END
   END FE_OFN286_n_29266

   PIN FE_OFN294_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.442 0.082 51.47 ;
      END
   END FE_OFN294_n_3069

   PIN FE_OFN331_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 55.922 0.163 55.95 ;
      END
   END FE_OFN331_n_4860

   PIN FE_OFN349_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.306 67.758 40.334 67.84 ;
      END
   END FE_OFN349_n_4860

   PIN FE_OFN37_n_17184
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 40.05 67.677 40.078 67.84 ;
      END
   END FE_OFN37_n_17184

   PIN FE_OFN404_n_28303
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 62.578 67.758 62.606 67.84 ;
      END
   END FE_OFN404_n_28303

   PIN FE_OFN68_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.438 27.89 99.52 27.918 ;
      END
   END FE_OFN68_n_27012

   PIN FE_OFN78_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 55.922 0.082 55.95 ;
      END
   END FE_OFN78_n_27012

   PIN FE_OFN7_n_28597
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.346 0.0 63.374 0.163 ;
      END
   END FE_OFN7_n_28597

   PIN FE_OFN95_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.762 0.0 43.79 0.082 ;
      END
   END FE_OFN95_n_27449

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 79.474 67.758 79.502 67.84 ;
      END
   END ispd_clk

   PIN n_1135
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.746 67.677 53.774 67.84 ;
      END
   END n_1135

   PIN n_11937
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.634 0.163 27.662 ;
      END
   END n_11937

   PIN n_12098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.754 0.163 24.782 ;
      END
   END n_12098

   PIN n_12562
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.73 0.163 39.758 ;
      END
   END n_12562

   PIN n_13053
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.618 0.163 13.646 ;
      END
   END n_13053

   PIN n_13876
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 55.666 0.163 55.694 ;
      END
   END n_13876

   PIN n_14512
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.602 0.163 39.63 ;
      END
   END n_14512

   PIN n_14515
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 46.578 0.163 46.606 ;
      END
   END n_14515

   PIN n_14997
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 73.202 67.677 73.23 67.84 ;
      END
   END n_14997

   PIN n_15183
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.738 67.677 26.766 67.84 ;
      END
   END n_15183

   PIN n_16917
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 42.162 0.163 42.19 ;
      END
   END n_16917

   PIN n_17248
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 60.466 0.163 60.494 ;
      END
   END n_17248

   PIN n_1774
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.378 67.677 59.406 67.84 ;
      END
   END n_1774

   PIN n_18484
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.002 0.163 62.03 ;
      END
   END n_18484

   PIN n_18834
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 41.842 0.163 41.87 ;
      END
   END n_18834

   PIN n_20042
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.866 0.163 18.894 ;
      END
   END n_20042

   PIN n_20287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.994 0.163 59.022 ;
      END
   END n_20287

   PIN n_21013
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 37.426 0.163 37.454 ;
      END
   END n_21013

   PIN n_21076
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.506 0.082 27.534 ;
      END
   END n_21076

   PIN n_21471
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.154 0.163 23.182 ;
      END
   END n_21471

   PIN n_21988
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 64.69 0.082 64.718 ;
      END
   END n_21988

   PIN n_22184
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.706 0.163 30.734 ;
      END
   END n_22184

   PIN n_22202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.626 0.163 32.654 ;
      END
   END n_22202

   PIN n_22681
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.258 0.163 62.286 ;
      END
   END n_22681

   PIN n_22758
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 27.826 0.163 27.854 ;
      END
   END n_22758

   PIN n_23465
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.762 0.163 27.79 ;
      END
   END n_23465

   PIN n_23509
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.602 67.677 79.63 67.84 ;
      END
   END n_23509

   PIN n_24114
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.698 0.163 27.726 ;
      END
   END n_24114

   PIN n_24126
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.418 0.163 18.446 ;
      END
   END n_24126

   PIN n_24135
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.498 0.163 32.526 ;
      END
   END n_24135

   PIN n_24421
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.33 67.677 89.358 67.84 ;
      END
   END n_24421

   PIN n_24716
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.802 0.163 18.83 ;
      END
   END n_24716

   PIN n_24799
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.274 67.677 84.302 67.84 ;
      END
   END n_24799

   PIN n_25130
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.146 67.677 84.174 67.84 ;
      END
   END n_25130

   PIN n_25150
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.546 0.163 18.574 ;
      END
   END n_25150

   PIN n_25188
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 53.554 99.52 53.582 ;
      END
   END n_25188

   PIN n_25502
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.978 67.677 85.006 67.84 ;
      END
   END n_25502

   PIN n_25659
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.626 0.163 8.654 ;
      END
   END n_25659

   PIN n_25660
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.69 0.163 8.718 ;
      END
   END n_25660

   PIN n_25661
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.818 0.163 8.846 ;
      END
   END n_25661

   PIN n_25854
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.202 0.163 17.23 ;
      END
   END n_25854

   PIN n_26081
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.626 67.677 80.654 67.84 ;
      END
   END n_26081

   PIN n_26139
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 51.314 99.52 51.342 ;
      END
   END n_26139

   PIN n_26416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 48.562 99.52 48.59 ;
      END
   END n_26416

   PIN n_26568
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.386 67.677 62.414 67.84 ;
      END
   END n_26568

   PIN n_26827
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 50.93 0.163 50.958 ;
      END
   END n_26827

   PIN n_26857
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 37.106 99.52 37.134 ;
      END
   END n_26857

   PIN n_27121
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 50.546 99.52 50.574 ;
      END
   END n_27121

   PIN n_27307
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 42.034 0.163 42.062 ;
      END
   END n_27307

   PIN n_27331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 60.53 0.163 60.558 ;
      END
   END n_27331

   PIN n_27332
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 97.586 67.677 97.614 67.84 ;
      END
   END n_27332

   PIN n_27415
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.362 67.677 69.39 67.84 ;
      END
   END n_27415

   PIN n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.922 67.758 55.95 67.84 ;
      END
   END n_27449

   PIN n_27488
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 76.786 67.677 76.814 67.84 ;
      END
   END n_27488

   PIN n_27709
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 73.906 0.0 73.934 0.082 ;
      END
   END n_27709

   PIN n_27914
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 50.802 0.163 50.83 ;
      END
   END n_27914

   PIN n_28602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 41.778 67.677 41.806 67.84 ;
      END
   END n_28602

   PIN n_28607
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 78.578 67.758 78.606 67.84 ;
      END
   END n_28607

   PIN n_29033
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.002 0.0 22.03 0.082 ;
      END
   END n_29033

   PIN n_29046
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 55.73 67.758 55.758 67.84 ;
      END
   END n_29046

   PIN n_29104
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 33.778 67.758 33.806 67.84 ;
      END
   END n_29104

   PIN n_29683
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.018 0.082 28.046 ;
      END
   END n_29683

   PIN n_29687
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 95.346 67.677 95.374 67.84 ;
      END
   END n_29687

   PIN n_29691
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.922 0.0 39.95 0.082 ;
      END
   END n_29691

   PIN n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.786 67.758 76.814 67.84 ;
      END
   END n_4280

   PIN n_4687
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 41.778 0.163 41.806 ;
      END
   END n_4687

   PIN n_4811
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.026 0.163 23.054 ;
      END
   END n_4811

   PIN n_5360
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.29 0.163 18.318 ;
      END
   END n_5360

   PIN n_5402
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 23.218 0.163 23.246 ;
      END
   END n_5402

   PIN n_5677
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.122 67.677 51.15 67.84 ;
      END
   END n_5677

   PIN n_5983
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 17.266 0.163 17.294 ;
      END
   END n_5983

   PIN n_6742
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.346 67.677 39.374 67.84 ;
      END
   END n_6742

   PIN n_6849
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 44.786 0.163 44.814 ;
      END
   END n_6849

   PIN n_7229
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.626 67.677 56.654 67.84 ;
      END
   END n_7229

   PIN n_7287
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.802 67.677 50.83 67.84 ;
      END
   END n_7287

   PIN n_7289
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.738 67.677 50.766 67.84 ;
      END
   END n_7289

   PIN n_7402
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.562 67.677 56.59 67.84 ;
      END
   END n_7402

   PIN n_7417
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.058 67.677 51.086 67.84 ;
      END
   END n_7417

   PIN n_8331
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.354 0.163 18.382 ;
      END
   END n_8331

   PIN n_8423
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.986 67.677 48.014 67.84 ;
      END
   END n_8423

   PIN n_8513
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.498 67.677 56.526 67.84 ;
      END
   END n_8513

   PIN n_8772
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.946 67.677 56.974 67.84 ;
      END
   END n_8772

   PIN n_8915
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 24.69 0.163 24.718 ;
      END
   END n_8915

   PIN n_9113
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.29 0.163 18.318 ;
      END
   END n_9113

   PIN n_9336
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 32.562 0.163 32.59 ;
      END
   END n_9336

   PIN n_9650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.482 0.163 18.51 ;
      END
   END n_9650

   PIN n_9936
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 18.738 0.163 18.766 ;
      END
   END n_9936

   PIN x_in_16_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 57.714 0.163 57.742 ;
      END
   END x_in_16_10

   PIN x_in_16_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 44.85 0.163 44.878 ;
      END
   END x_in_16_11

   PIN x_in_16_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 33.394 0.163 33.422 ;
      END
   END x_in_16_12

   PIN x_in_16_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 19.314 0.163 19.342 ;
      END
   END x_in_16_13

   PIN x_in_16_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.994 0.163 19.022 ;
      END
   END x_in_16_14

   PIN x_in_16_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.426 0.163 13.454 ;
      END
   END x_in_16_15

   PIN x_in_16_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 4.914 67.677 4.942 67.84 ;
      END
   END x_in_16_3

   PIN x_in_16_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 65.202 0.163 65.23 ;
      END
   END x_in_16_4

   PIN x_in_16_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 53.682 0.163 53.71 ;
      END
   END x_in_16_5

   PIN x_in_16_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 14.258 67.677 14.286 67.84 ;
      END
   END x_in_16_6

   PIN x_in_16_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 56.05 0.163 56.078 ;
      END
   END x_in_16_7

   PIN x_in_17_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 8.754 0.163 8.782 ;
      END
   END x_in_17_15

   PIN x_in_17_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.89 0.163 27.918 ;
      END
   END x_in_17_2

   PIN x_in_17_3
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 45.17 0.082 45.198 ;
      END
   END x_in_17_3

   PIN x_in_17_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 46.258 0.082 46.286 ;
      END
   END x_in_17_4

   PIN x_in_17_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 27.698 0.082 27.726 ;
      END
   END x_in_17_5

   PIN x_in_17_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 31.282 0.082 31.31 ;
      END
   END x_in_17_6

   PIN x_in_17_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 21.81 0.082 21.838 ;
      END
   END x_in_17_7

   PIN x_in_17_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 18.418 0.082 18.446 ;
      END
   END x_in_17_8

   PIN x_in_26_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.226 67.677 82.254 67.84 ;
      END
   END x_in_26_10

   PIN x_in_26_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 62.194 0.163 62.222 ;
      END
   END x_in_26_11

   PIN x_in_26_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 99.357 46.514 99.52 46.542 ;
      END
   END x_in_26_12

   PIN x_in_26_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 36.338 0.163 36.366 ;
      END
   END x_in_26_13

   PIN x_in_26_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.722 0.163 36.75 ;
      END
   END x_in_26_14

   PIN x_in_26_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 62.13 0.163 62.158 ;
      END
   END x_in_26_15

   PIN x_in_27_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.866 67.677 50.894 67.84 ;
      END
   END x_in_27_10

   PIN x_in_27_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 50.866 67.758 50.894 67.84 ;
      END
   END x_in_27_11

   PIN x_in_27_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.506 67.677 59.534 67.84 ;
      END
   END x_in_27_12

   PIN x_in_27_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.474 67.677 63.502 67.84 ;
      END
   END x_in_27_13

   PIN x_in_27_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.442 67.677 59.47 67.84 ;
      END
   END x_in_27_14

   PIN x_in_27_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 58.226 67.677 58.254 67.84 ;
      END
   END x_in_27_15

   PIN x_in_27_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 53.81 67.677 53.838 67.84 ;
      END
   END x_in_27_9

   PIN x_out_22_21
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.042 67.677 45.07 67.84 ;
      END
   END x_out_22_21

   PIN x_out_22_22
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 88.37 67.677 88.398 67.84 ;
      END
   END x_out_22_22

   PIN x_out_2_31
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.466 67.677 28.494 67.84 ;
      END
   END x_out_2_31

   PIN x_out_34_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 48.818 0.163 48.846 ;
      END
   END x_out_34_12

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 99.52 67.84 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 99.52 67.84 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 99.52 67.84 ;
      LAYER V1 ;
         RECT 0.0 0.0 99.52 67.84 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 99.52 67.84 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 99.52 67.84 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 99.52 67.84 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 99.52 67.84 ;
      LAYER M1 ;
         RECT 0.0 0.0 99.52 67.84 ;
   END
END h4_mgc_fft_a

MACRO h3_mgc_fft_a
   CLASS BLOCK ;
   FOREIGN h3 ;
   ORIGIN 0 0 ;
   SIZE 222.976 BY 55.04 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1143_n_27012
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 175.026 0.0 175.054 0.082 ;
      END
   END FE_OFN1143_n_27012

   PIN FE_OFN1193_n_12908
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.01 0.0 129.038 0.163 ;
      END
   END FE_OFN1193_n_12908

   PIN FE_OFN612_n_5698
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.314 54.877 51.342 55.04 ;
      END
   END FE_OFN612_n_5698

   PIN FE_OFN734_n_22952
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.77 0.163 30.798 ;
      END
   END FE_OFN734_n_22952

   PIN FE_OFN750_n_20252
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.674 0.0 42.702 0.163 ;
      END
   END FE_OFN750_n_20252

   PIN n_10335
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.81 0.0 13.838 0.163 ;
      END
   END n_10335

   PIN n_10432
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 124.658 0.0 124.686 0.163 ;
      END
   END n_10432

   PIN n_11256
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.482 54.877 34.51 55.04 ;
      END
   END n_11256

   PIN n_11262
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 13.554 222.976 13.582 ;
      END
   END n_11262

   PIN n_11285
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.794 54.877 39.822 55.04 ;
      END
   END n_11285

   PIN n_11526
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 221.17 0.0 221.198 0.163 ;
      END
   END n_11526

   PIN n_12365
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.514 0.0 126.542 0.163 ;
      END
   END n_12365

   PIN n_12646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 27.506 222.976 27.534 ;
      END
   END n_12646

   PIN n_13045
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.666 54.877 39.694 55.04 ;
      END
   END n_13045

   PIN n_13066
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 8.05 0.0 8.078 0.163 ;
      END
   END n_13066

   PIN n_13175
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.362 0.0 5.39 0.163 ;
      END
   END n_13175

   PIN n_13229
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.186 54.877 51.214 55.04 ;
      END
   END n_13229

   PIN n_13260
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.946 54.877 56.974 55.04 ;
      END
   END n_13260

   PIN n_1333
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.874 54.877 13.902 55.04 ;
      END
   END n_1333

   PIN n_13379
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 212.53 0.0 212.558 0.163 ;
      END
   END n_13379

   PIN n_13564
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 154.034 0.0 154.062 0.163 ;
      END
   END n_13564

   PIN n_13965
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.186 0.0 123.214 0.163 ;
      END
   END n_13965

   PIN n_14028
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 13.618 222.976 13.646 ;
      END
   END n_14028

   PIN n_14346
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.002 54.877 38.03 55.04 ;
      END
   END n_14346

   PIN n_14354
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 139.698 0.0 139.726 0.163 ;
      END
   END n_14354

   PIN n_14355
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 140.53 0.0 140.558 0.163 ;
      END
   END n_14355

   PIN n_14407
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 3.314 0.0 3.342 0.163 ;
      END
   END n_14407

   PIN n_14580
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.85 54.877 180.878 55.04 ;
      END
   END n_14580

   PIN n_14926
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 22.194 222.976 22.222 ;
      END
   END n_14926

   PIN n_14927
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 30.834 222.976 30.862 ;
      END
   END n_14927

   PIN n_15065
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 16.562 222.976 16.59 ;
      END
   END n_15065

   PIN n_15131
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.89 54.877 35.918 55.04 ;
      END
   END n_15131

   PIN n_15879
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.234 0.0 5.262 0.163 ;
      END
   END n_15879

   PIN n_15880
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.354 0.0 2.382 0.163 ;
      END
   END n_15880

   PIN n_15991
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 175.09 54.877 175.118 55.04 ;
      END
   END n_15991

   PIN n_16350
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.29 0.0 146.318 0.163 ;
      END
   END n_16350

   PIN n_16586
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 2.29 0.0 2.318 0.163 ;
      END
   END n_16586

   PIN n_16635
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 175.09 54.877 175.118 55.04 ;
      END
   END n_16635

   PIN n_16639
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.026 54.877 135.054 55.04 ;
      END
   END n_16639

   PIN n_16640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.898 54.877 134.926 55.04 ;
      END
   END n_16640

   PIN n_16886
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.962 54.877 134.99 55.04 ;
      END
   END n_16886

   PIN n_17035
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.194 0.163 22.222 ;
      END
   END n_17035

   PIN n_17253
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 45.234 222.976 45.262 ;
      END
   END n_17253

   PIN n_17495
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.89 54.877 131.918 55.04 ;
      END
   END n_17495

   PIN n_18101
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.018 0.163 4.046 ;
      END
   END n_18101

   PIN n_18104
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 39.474 222.976 39.502 ;
      END
   END n_18104

   PIN n_18396
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.066 0.0 126.094 0.163 ;
      END
   END n_18396

   PIN n_18435
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 45.298 222.976 45.326 ;
      END
   END n_18435

   PIN n_18488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.146 0.163 4.174 ;
      END
   END n_18488

   PIN n_18650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.498 0.0 8.526 0.163 ;
      END
   END n_18650

   PIN n_18683
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.45 0.0 126.478 0.163 ;
      END
   END n_18683

   PIN n_18728
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 209.65 54.877 209.678 55.04 ;
      END
   END n_18728

   PIN n_18812
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.562 0.163 16.59 ;
      END
   END n_18812

   PIN n_18882
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.506 0.163 27.534 ;
      END
   END n_18882

   PIN n_19039
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.906 54.877 33.934 55.04 ;
      END
   END n_19039

   PIN n_19298
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 10.098 0.0 10.126 0.163 ;
      END
   END n_19298

   PIN n_19968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.21 0.0 28.238 0.163 ;
      END
   END n_19968

   PIN n_20250
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.146 0.0 20.174 0.163 ;
      END
   END n_20250

   PIN n_20474
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 116.274 0.0 116.302 0.163 ;
      END
   END n_20474

   PIN n_20562
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.898 0.0 38.926 0.163 ;
      END
   END n_20562

   PIN n_20792
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.122 0.163 3.15 ;
      END
   END n_20792

   PIN n_20875
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 171.826 0.0 171.854 0.163 ;
      END
   END n_20875

   PIN n_21178
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.73 54.877 39.758 55.04 ;
      END
   END n_21178

   PIN n_21295
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.634 0.163 19.662 ;
      END
   END n_21295

   PIN n_21341
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.578 0.0 22.606 0.163 ;
      END
   END n_21341

   PIN n_21463
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.634 0.0 67.662 0.163 ;
      END
   END n_21463

   PIN n_21562
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 35.122 222.976 35.15 ;
      END
   END n_21562

   PIN n_21991
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.514 54.877 166.542 55.04 ;
      END
   END n_21991

   PIN n_2220
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.01 0.0 201.038 0.163 ;
      END
   END n_2220

   PIN n_23291
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.274 0.0 44.302 0.082 ;
      END
   END n_23291

   PIN n_2342
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 192.37 0.0 192.398 0.163 ;
      END
   END n_2342

   PIN n_24279
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.89 0.163 3.918 ;
      END
   END n_24279

   PIN n_24915
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.546 0.0 82.574 0.163 ;
      END
   END n_24915

   PIN n_25379
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.33 0.0 25.358 0.163 ;
      END
   END n_25379

   PIN n_25402
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.266 0.0 25.294 0.163 ;
      END
   END n_25402

   PIN n_25645
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.914 0.0 52.942 0.163 ;
      END
   END n_25645

   PIN n_27432
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.914 0.0 36.942 0.163 ;
      END
   END n_27432

   PIN n_276
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.922 0.0 39.95 0.163 ;
      END
   END n_276

   PIN n_27650
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 84.658 0.0 84.686 0.163 ;
      END
   END n_27650

   PIN n_27750
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 30.834 0.163 30.862 ;
      END
   END n_27750

   PIN n_28369
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.354 0.0 82.382 0.163 ;
      END
   END n_28369

   PIN n_3620
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 52.85 54.877 52.878 55.04 ;
      END
   END n_3620

   PIN n_3621
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.586 54.877 57.614 55.04 ;
      END
   END n_3621

   PIN n_3811
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 192.434 0.0 192.462 0.163 ;
      END
   END n_3811

   PIN n_3847
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 188.914 0.0 188.942 0.163 ;
      END
   END n_3847

   PIN n_4099
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 122.866 0.0 122.894 0.163 ;
      END
   END n_4099

   PIN n_4578
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.874 0.0 13.902 0.163 ;
      END
   END n_4578

   PIN n_4928
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.666 0.0 119.694 0.163 ;
      END
   END n_4928

   PIN n_5156
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.698 0.0 11.726 0.163 ;
      END
   END n_5156

   PIN n_5158
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.866 0.0 10.894 0.163 ;
      END
   END n_5158

   PIN n_5537
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.322 54.877 38.35 55.04 ;
      END
   END n_5537

   PIN n_5556
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.378 54.877 51.406 55.04 ;
      END
   END n_5556

   PIN n_5557
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.25 54.877 51.278 55.04 ;
      END
   END n_5557

   PIN n_5601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.674 0.0 186.702 0.163 ;
      END
   END n_5601

   PIN n_5602
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 186.61 0.0 186.638 0.163 ;
      END
   END n_5602

   PIN n_5637
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 198.13 0.0 198.158 0.163 ;
      END
   END n_5637

   PIN n_5689
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.41 0.0 215.438 0.163 ;
      END
   END n_5689

   PIN n_5794
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.642 54.877 134.67 55.04 ;
      END
   END n_5794

   PIN n_5845
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.898 54.877 54.926 55.04 ;
      END
   END n_5845

   PIN n_5928
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.066 54.877 54.094 55.04 ;
      END
   END n_5928

   PIN n_6420
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 203.89 0.0 203.918 0.163 ;
      END
   END n_6420

   PIN n_6538
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.146 54.877 60.174 55.04 ;
      END
   END n_6538

   PIN n_6631
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 123.25 0.0 123.278 0.163 ;
      END
   END n_6631

   PIN n_6646
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 134.706 54.877 134.734 55.04 ;
      END
   END n_6646

   PIN n_7384
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 8.05 0.0 8.078 0.163 ;
      END
   END n_7384

   PIN n_8420
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 181.234 0.0 181.262 0.163 ;
      END
   END n_8420

   PIN n_9616
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 206.834 0.0 206.862 0.163 ;
      END
   END n_9616

   PIN n_9619
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 109.106 0.0 109.134 0.163 ;
      END
   END n_9619

   PIN n_9640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.858 54.877 39.886 55.04 ;
      END
   END n_9640

   PIN n_9641
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.794 54.877 39.822 55.04 ;
      END
   END n_9641

   PIN n_9644
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.434 54.877 48.462 55.04 ;
      END
   END n_9644

   PIN n_9838
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 19.634 222.976 19.662 ;
      END
   END n_9838

   PIN n_9937
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.986 54.877 80.014 55.04 ;
      END
   END n_9937

   PIN n_999
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.442 0.163 43.47 ;
      END
   END n_999

   PIN x_out_12_27
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 183.73 0.0 183.758 0.163 ;
      END
   END x_out_12_27

   PIN x_out_12_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.37 54.877 120.398 55.04 ;
      END
   END x_out_12_28

   PIN x_out_12_31
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 180.914 0.0 180.942 0.163 ;
      END
   END x_out_12_31

   PIN x_out_17_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.682 0.163 13.71 ;
      END
   END x_out_17_24

   PIN x_out_17_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.714 0.0 65.742 0.163 ;
      END
   END x_out_17_7

   PIN x_out_17_8
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 13.49 0.163 13.518 ;
      END
   END x_out_17_8

   PIN x_out_18_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 48.05 0.163 48.078 ;
      END
   END x_out_18_1

   PIN x_out_18_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 28.274 0.0 28.302 0.163 ;
      END
   END x_out_18_12

   PIN x_out_1_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.05 0.0 88.078 0.163 ;
      END
   END x_out_1_11

   PIN x_out_30_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 180.85 0.0 180.878 0.163 ;
      END
   END x_out_30_3

   PIN x_out_30_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 166.45 0.0 166.478 0.163 ;
      END
   END x_out_30_4

   PIN x_out_33_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.514 0.0 22.542 0.163 ;
      END
   END x_out_33_10

   PIN x_out_33_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.45 0.0 22.478 0.163 ;
      END
   END x_out_33_12

   PIN x_out_42_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 80.114 0.0 80.142 0.163 ;
      END
   END x_out_42_24

   PIN x_out_44_23
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 152.562 0.0 152.59 0.163 ;
      END
   END x_out_44_23

   PIN x_out_44_26
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 172.146 0.0 172.174 0.163 ;
      END
   END x_out_44_26

   PIN x_out_49_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 10.546 0.163 10.574 ;
      END
   END x_out_49_10

   PIN x_out_49_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 4.914 0.163 4.942 ;
      END
   END x_out_49_24

   PIN x_out_49_32
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.034 0.0 34.062 0.163 ;
      END
   END x_out_49_32

   PIN x_out_62_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 200.946 0.0 200.974 0.163 ;
      END
   END x_out_62_11

   PIN FE_OFN1123_rst
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 95.026 0.0 95.054 0.082 ;
      END
   END FE_OFN1123_rst

   PIN FE_OFN1124_rst
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.746 0.0 85.774 0.082 ;
      END
   END FE_OFN1124_rst

   PIN FE_OFN116_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 186.61 0.0 186.638 0.082 ;
      END
   END FE_OFN116_n_27449

   PIN FE_OFN1181_rst
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 192.69 54.958 192.718 55.04 ;
      END
   END FE_OFN1181_rst

   PIN FE_OFN129_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 169.33 0.0 169.358 0.082 ;
      END
   END FE_OFN129_n_27449

   PIN FE_OFN131_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 35.378 0.082 35.406 ;
      END
   END FE_OFN131_n_27449

   PIN FE_OFN139_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 38.066 0.0 38.094 0.082 ;
      END
   END FE_OFN139_n_27449

   PIN FE_OFN173_n_22948
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.61 0.0 42.638 0.163 ;
      END
   END FE_OFN173_n_22948

   PIN FE_OFN199_n_29637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 175.154 0.0 175.182 0.163 ;
      END
   END FE_OFN199_n_29637

   PIN FE_OFN206_n_28771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 170.162 54.877 170.19 55.04 ;
      END
   END FE_OFN206_n_28771

   PIN FE_OFN235_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 192.498 54.958 192.526 55.04 ;
      END
   END FE_OFN235_n_4162

   PIN FE_OFN23_n_26609
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 90.546 0.0 90.574 0.163 ;
      END
   END FE_OFN23_n_26609

   PIN FE_OFN244_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 37.874 0.0 37.902 0.082 ;
      END
   END FE_OFN244_n_4162

   PIN FE_OFN254_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 65.842 0.0 65.87 0.082 ;
      END
   END FE_OFN254_n_4280

   PIN FE_OFN266_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 150.386 54.958 150.414 55.04 ;
      END
   END FE_OFN266_n_4280

   PIN FE_OFN280_n_16656
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 103.09 54.877 103.118 55.04 ;
      END
   END FE_OFN280_n_16656

   PIN FE_OFN296_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 82.29 54.958 82.318 55.04 ;
      END
   END FE_OFN296_n_3069

   PIN FE_OFN310_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 169.266 54.958 169.294 55.04 ;
      END
   END FE_OFN310_n_3069

   PIN FE_OFN313_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 34.162 0.0 34.19 0.082 ;
      END
   END FE_OFN313_n_3069

   PIN FE_OFN335_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 175.346 0.0 175.374 0.082 ;
      END
   END FE_OFN335_n_4860

   PIN FE_OFN361_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 80.626 54.958 80.654 55.04 ;
      END
   END FE_OFN361_n_4860

   PIN FE_OFN3_n_28682
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.858 0.0 31.886 0.163 ;
      END
   END FE_OFN3_n_28682

   PIN FE_OFN4_n_28682
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 182.258 0.0 182.286 0.163 ;
      END
   END FE_OFN4_n_28682

   PIN FE_OFN553_n_9468
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 149.17 0.0 149.198 0.163 ;
      END
   END FE_OFN553_n_9468

   PIN FE_OFN56_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 195.314 0.0 195.342 0.082 ;
      END
   END FE_OFN56_n_27012

   PIN FE_OFN63_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 165.618 0.0 165.646 0.082 ;
      END
   END FE_OFN63_n_27012

   PIN FE_OFN695_n_19853
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 48.114 222.976 48.142 ;
      END
   END FE_OFN695_n_19853

   PIN FE_OFN733_n_22952
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.154 0.0 31.182 0.163 ;
      END
   END FE_OFN733_n_22952

   PIN FE_OFN80_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 39.73 0.0 39.758 0.082 ;
      END
   END FE_OFN80_n_27012

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 178.226 0.0 178.254 0.082 ;
      END
   END ispd_clk

   PIN n_10089
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 176.434 0.0 176.462 0.163 ;
      END
   END n_10089

   PIN n_10416
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 35.314 222.976 35.342 ;
      END
   END n_10416

   PIN n_10590
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.13 54.877 38.158 55.04 ;
      END
   END n_10590

   PIN n_10591
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.842 54.877 33.87 55.04 ;
      END
   END n_10591

   PIN n_10729
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 107.25 0.0 107.278 0.163 ;
      END
   END n_10729

   PIN n_10751
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.938 0.0 13.966 0.163 ;
      END
   END n_10751

   PIN n_11036
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.17 0.0 5.198 0.163 ;
      END
   END n_11036

   PIN n_11157
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.618 0.0 13.646 0.163 ;
      END
   END n_11157

   PIN n_11245
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.522 0.0 25.55 0.163 ;
      END
   END n_11245

   PIN n_11246
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.386 0.0 22.414 0.163 ;
      END
   END n_11246

   PIN n_11255
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.546 54.877 34.574 55.04 ;
      END
   END n_11255

   PIN n_11257
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.962 54.877 30.99 55.04 ;
      END
   END n_11257

   PIN n_11258
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.37 54.877 48.398 55.04 ;
      END
   END n_11258

   PIN n_11261
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 27.57 222.976 27.598 ;
      END
   END n_11261

   PIN n_11288
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.634 0.0 19.662 0.163 ;
      END
   END n_11288

   PIN n_11289
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.57 0.0 19.598 0.163 ;
      END
   END n_11289

   PIN n_11700
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 155.25 0.0 155.278 0.163 ;
      END
   END n_11700

   PIN n_11930
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.938 0.0 157.966 0.163 ;
      END
   END n_11930

   PIN n_12647
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 27.442 222.976 27.47 ;
      END
   END n_12647

   PIN n_12770
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.93 0.0 18.958 0.163 ;
      END
   END n_12770

   PIN n_12860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.242 0.0 160.27 0.163 ;
      END
   END n_12860

   PIN n_12861
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.05 0.0 160.078 0.163 ;
      END
   END n_12861

   PIN n_13489
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 160.178 0.0 160.206 0.163 ;
      END
   END n_13489

   PIN n_13775
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 169.33 0.0 169.358 0.163 ;
      END
   END n_13775

   PIN n_15151
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 1.266 0.0 1.294 0.163 ;
      END
   END n_15151

   PIN n_15466
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 222.813 45.234 222.976 45.262 ;
      END
   END n_15466

   PIN n_15467
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 43.442 222.976 43.47 ;
      END
   END n_15467

   PIN n_15726
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 50.994 222.976 51.022 ;
      END
   END n_15726

   PIN n_15952
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.298 0.0 5.326 0.163 ;
      END
   END n_15952

   PIN n_16194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 45.17 222.976 45.198 ;
      END
   END n_16194

   PIN n_16346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 173.81 54.877 173.838 55.04 ;
      END
   END n_16346

   PIN n_16852
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.29 0.0 2.318 0.163 ;
      END
   END n_16852

   PIN n_17198
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 81.01 0.0 81.038 0.163 ;
      END
   END n_17198

   PIN n_17337
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 7.794 0.163 7.822 ;
      END
   END n_17337

   PIN n_17343
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 48.242 222.976 48.27 ;
      END
   END n_17343

   PIN n_17394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 22.13 0.163 22.158 ;
      END
   END n_17394

   PIN n_17493
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 180.914 54.877 180.942 55.04 ;
      END
   END n_17493

   PIN n_17810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.93 54.877 130.958 55.04 ;
      END
   END n_17810

   PIN n_17907
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 4.082 0.163 4.11 ;
      END
   END n_17907

   PIN n_18098
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 126.45 54.877 126.478 55.04 ;
      END
   END n_18098

   PIN n_18350
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.442 0.0 19.47 0.163 ;
      END
   END n_18350

   PIN n_18487
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 3.954 0.163 3.982 ;
      END
   END n_18487

   PIN n_18727
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 210.226 54.877 210.254 55.04 ;
      END
   END n_18727

   PIN n_1878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 166.45 54.877 166.478 55.04 ;
      END
   END n_1878

   PIN n_18914
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.034 0.0 10.062 0.163 ;
      END
   END n_18914

   PIN n_18915
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.226 0.0 10.254 0.163 ;
      END
   END n_18915

   PIN n_19090
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 48.178 222.976 48.206 ;
      END
   END n_19090

   PIN n_19923
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.802 0.163 10.83 ;
      END
   END n_19923

   PIN n_20095
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.97 54.877 33.998 55.04 ;
      END
   END n_20095

   PIN n_20160
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 222.813 45.298 222.976 45.326 ;
      END
   END n_20160

   PIN n_20293
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 64.498 0.0 64.526 0.163 ;
      END
   END n_20293

   PIN n_20322
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 5.17 54.877 5.198 55.04 ;
      END
   END n_20322

   PIN n_20561
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.962 0.0 38.99 0.163 ;
      END
   END n_20561

   PIN n_20563
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 38.77 0.0 38.798 0.163 ;
      END
   END n_20563

   PIN n_20717
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.89 0.0 59.918 0.163 ;
      END
   END n_20717

   PIN n_20876
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 170.546 0.0 170.574 0.163 ;
      END
   END n_20876

   PIN n_20978
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.506 0.0 19.534 0.163 ;
      END
   END n_20978

   PIN n_21000
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.09 0.0 31.118 0.163 ;
      END
   END n_21000

   PIN n_22275
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.026 0.0 31.054 0.163 ;
      END
   END n_22275

   PIN n_24278
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 3.89 0.163 3.918 ;
      END
   END n_24278

   PIN n_24691
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.25 0.0 27.278 0.163 ;
      END
   END n_24691

   PIN n_24916
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.33 0.0 25.358 0.163 ;
      END
   END n_24916

   PIN n_25378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.202 0.0 25.23 0.163 ;
      END
   END n_25378

   PIN n_25680
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 150.514 54.958 150.542 55.04 ;
      END
   END n_25680

   PIN n_25987
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 85.618 0.0 85.646 0.163 ;
      END
   END n_25987

   PIN n_26637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 2.418 0.0 2.446 0.163 ;
      END
   END n_26637

   PIN n_2673
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 135.538 0.0 135.566 0.163 ;
      END
   END n_2673

   PIN n_2696
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 205.298 0.0 205.326 0.163 ;
      END
   END n_2696

   PIN n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 206.77 54.958 206.798 55.04 ;
      END
   END n_27012

   PIN n_27270
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.97 0.0 33.998 0.163 ;
      END
   END n_27270

   PIN n_27933
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 195.122 0.0 195.15 0.082 ;
      END
   END n_27933

   PIN n_28094
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.474 0.163 39.502 ;
      END
   END n_28094

   PIN n_28101
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 45.234 0.163 45.262 ;
      END
   END n_28101

   PIN n_28102
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.298 0.163 45.326 ;
      END
   END n_28102

   PIN n_28263
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.234 0.163 45.262 ;
      END
   END n_28263

   PIN n_28319
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.85 0.0 36.878 0.163 ;
      END
   END n_28319

   PIN n_28325
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.73 0.0 31.758 0.163 ;
      END
   END n_28325

   PIN n_28330
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 222.813 30.77 222.976 30.798 ;
      END
   END n_28330

   PIN n_2834
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.306 0.0 120.334 0.163 ;
      END
   END n_2834

   PIN n_28362
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.482 54.877 82.51 55.04 ;
      END
   END n_28362

   PIN n_29100
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.81 54.877 13.838 55.04 ;
      END
   END n_29100

   PIN n_3020
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 45.49 54.877 45.518 55.04 ;
      END
   END n_3020

   PIN n_3082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.77 54.877 62.798 55.04 ;
      END
   END n_3082

   PIN n_3781
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.674 54.877 42.702 55.04 ;
      END
   END n_3781

   PIN n_3853
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.026 0.0 119.054 0.163 ;
      END
   END n_3853

   PIN n_4057
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 67.378 54.877 67.406 55.04 ;
      END
   END n_4057

   PIN n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 150.834 54.958 150.862 55.04 ;
      END
   END n_4162

   PIN n_4270
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 44.338 54.958 44.366 55.04 ;
      END
   END n_4270

   PIN n_4400
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 42.61 54.877 42.638 55.04 ;
      END
   END n_4400

   PIN n_4454
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.626 0.0 160.654 0.163 ;
      END
   END n_4454

   PIN n_4577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.746 0.0 13.774 0.163 ;
      END
   END n_4577

   PIN n_4890
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 118.834 0.0 118.862 0.163 ;
      END
   END n_4890

   PIN n_4929
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 119.73 0.0 119.758 0.163 ;
      END
   END n_4929

   PIN n_5157
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.13 0.0 22.158 0.163 ;
      END
   END n_5157

   PIN n_5243
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.122 54.877 51.15 55.04 ;
      END
   END n_5243

   PIN n_5264
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 155.442 0.0 155.47 0.163 ;
      END
   END n_5264

   PIN n_5283
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 218.29 0.0 218.318 0.163 ;
      END
   END n_5283

   PIN n_5338
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.49 0.0 117.518 0.163 ;
      END
   END n_5338

   PIN n_5487
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 47.794 54.877 47.822 55.04 ;
      END
   END n_5487

   PIN n_5539
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.938 54.877 29.966 55.04 ;
      END
   END n_5539

   PIN n_5554
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 45.426 54.877 45.454 55.04 ;
      END
   END n_5554

   PIN n_5664
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.066 54.877 30.094 55.04 ;
      END
   END n_5664

   PIN n_5925
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 120.242 0.0 120.27 0.163 ;
      END
   END n_5925

   PIN n_5926
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 117.426 0.0 117.454 0.163 ;
      END
   END n_5926

   PIN n_6258
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.602 54.877 39.63 55.04 ;
      END
   END n_6258

   PIN n_6285
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 117.49 0.0 117.518 0.163 ;
      END
   END n_6285

   PIN n_6311
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 201.778 0.0 201.806 0.163 ;
      END
   END n_6311

   PIN n_7765
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.114 54.958 48.142 55.04 ;
      END
   END n_7765

   PIN n_7796
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.002 54.877 30.03 55.04 ;
      END
   END n_7796

   PIN n_7797
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.474 54.877 23.502 55.04 ;
      END
   END n_7797

   PIN n_7802
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.306 54.877 48.334 55.04 ;
      END
   END n_7802

   PIN n_7810
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 200.946 0.0 200.974 0.163 ;
      END
   END n_7810

   PIN n_7823
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.73 54.877 39.758 55.04 ;
      END
   END n_7823

   PIN n_8345
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 11.25 0.0 11.278 0.163 ;
      END
   END n_8345

   PIN n_8346
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 10.802 0.0 10.83 0.163 ;
      END
   END n_8346

   PIN n_8489
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.026 0.0 23.054 0.163 ;
      END
   END n_8489

   PIN n_8490
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.562 0.0 16.59 0.163 ;
      END
   END n_8490

   PIN n_8919
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 14.002 0.0 14.03 0.163 ;
      END
   END n_8919

   PIN n_8920
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.626 0.0 16.654 0.163 ;
      END
   END n_8920

   PIN n_9440
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 215.474 0.0 215.502 0.163 ;
      END
   END n_9440

   PIN n_9482
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 157.81 0.0 157.838 0.163 ;
      END
   END n_9482

   PIN n_9617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 194.482 0.0 194.51 0.163 ;
      END
   END n_9617

   PIN n_9637
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 29.746 54.877 29.774 55.04 ;
      END
   END n_9637

   PIN n_9645
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.242 54.877 48.27 55.04 ;
      END
   END n_9645

   PIN n_9662
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.922 0.0 15.95 0.163 ;
      END
   END n_9662

   PIN n_9663
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 15.858 0.0 15.886 0.163 ;
      END
   END n_9663

   PIN n_9664
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.682 0.0 13.71 0.163 ;
      END
   END n_9664

   PIN n_9737
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.57 0.0 19.598 0.163 ;
      END
   END n_9737

   PIN n_9961
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.818 0.0 16.846 0.163 ;
      END
   END n_9961

   PIN x_in_13_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 130.098 0.0 130.126 0.163 ;
      END
   END x_in_13_10

   PIN x_in_13_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 135.474 0.0 135.502 0.082 ;
      END
   END x_in_13_11

   PIN x_in_13_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 123.25 0.0 123.278 0.163 ;
      END
   END x_in_13_12

   PIN x_in_13_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 131.954 0.0 131.982 0.163 ;
      END
   END x_in_13_13

   PIN x_in_13_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 129.074 0.0 129.102 0.163 ;
      END
   END x_in_13_14

   PIN x_in_13_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 160.754 0.0 160.782 0.163 ;
      END
   END x_in_13_9

   PIN x_in_19_10
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.026 54.958 31.054 55.04 ;
      END
   END x_in_19_10

   PIN x_in_19_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.37 54.958 48.398 55.04 ;
      END
   END x_in_19_11

   PIN x_in_19_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 54.322 54.958 54.35 55.04 ;
      END
   END x_in_19_12

   PIN x_in_19_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 54.066 54.958 54.094 55.04 ;
      END
   END x_in_19_13

   PIN x_in_19_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.714 54.877 57.742 55.04 ;
      END
   END x_in_19_14

   PIN x_in_19_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 54.194 54.877 54.222 55.04 ;
      END
   END x_in_19_15

   PIN x_in_19_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.826 54.958 43.854 55.04 ;
      END
   END x_in_19_9

   PIN x_in_30_2
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 166.514 0.0 166.542 0.163 ;
      END
   END x_in_30_2

   PIN x_in_34_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 13.554 0.163 13.582 ;
      END
   END x_in_34_7

   PIN x_in_35_1
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 16.69 0.0 16.718 0.082 ;
      END
   END x_in_35_1

   PIN x_in_51_11
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 198.194 0.0 198.222 0.082 ;
      END
   END x_in_51_11

   PIN x_in_51_12
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 206.642 0.0 206.67 0.082 ;
      END
   END x_in_51_12

   PIN x_in_51_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 201.074 0.0 201.102 0.163 ;
      END
   END x_in_51_13

   PIN x_in_51_14
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 198.066 0.0 198.094 0.163 ;
      END
   END x_in_51_14

   PIN x_in_51_15
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 206.77 0.0 206.798 0.163 ;
      END
   END x_in_51_15

   PIN x_out_12_26
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 146.354 0.0 146.382 0.163 ;
      END
   END x_out_12_26

   PIN x_out_49_30
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 82.738 0.0 82.766 0.163 ;
      END
   END x_out_49_30

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 222.976 55.04 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 222.976 55.04 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 222.976 55.04 ;
      LAYER V1 ;
         RECT 0.0 0.0 222.976 55.04 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 222.976 55.04 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 222.976 55.04 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 222.976 55.04 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 222.976 55.04 ;
      LAYER M1 ;
         RECT 0.0 0.0 222.976 55.04 ;
   END
END h3_mgc_fft_a

MACRO h2_mgc_fft_a
   CLASS BLOCK ;
   FOREIGN h2 ;
   ORIGIN 0 0 ;
   SIZE 106.432 BY 81.28 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN953_n_13421
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 13.618 81.117 13.646 81.28 ;
      END
   END FE_OFN953_n_13421

   PIN n_10046
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 31.282 0.163 31.31 ;
      END
   END n_10046

   PIN n_10214
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 11.122 0.163 11.15 ;
      END
   END n_10214

   PIN n_1203
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.778 81.117 25.806 81.28 ;
      END
   END n_1203

   PIN n_12798
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.914 0.163 36.942 ;
      END
   END n_12798

   PIN n_13206
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.554 0.163 45.582 ;
      END
   END n_13206

   PIN n_13818
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.474 81.117 31.502 81.28 ;
      END
   END n_13818

   PIN n_14891
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 31.602 81.117 31.63 81.28 ;
      END
   END n_14891

   PIN n_15558
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 15.474 81.117 15.502 81.28 ;
      END
   END n_15558

   PIN n_19720
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 19.506 81.117 19.534 81.28 ;
      END
   END n_19720

   PIN n_21108
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.922 81.117 23.95 81.28 ;
      END
   END n_21108

   PIN n_21121
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.522 81.117 17.55 81.28 ;
      END
   END n_21121

   PIN n_23262
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.146 81.117 20.174 81.28 ;
      END
   END n_23262

   PIN n_23263
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.018 81.117 20.046 81.28 ;
      END
   END n_23263

   PIN n_23336
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 26.098 81.117 26.126 81.28 ;
      END
   END n_23336

   PIN n_24991
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 20.082 81.117 20.11 81.28 ;
      END
   END n_24991

   PIN n_25847
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.418 81.117 34.446 81.28 ;
      END
   END n_25847

   PIN n_26581
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.41 81.117 31.438 81.28 ;
      END
   END n_26581

   PIN n_26926
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.986 81.117 32.014 81.28 ;
      END
   END n_26926

   PIN n_29040
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 59.954 0.163 59.982 ;
      END
   END n_29040

   PIN n_29135
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.33 81.117 33.358 81.28 ;
      END
   END n_29135

   PIN n_4730
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.442 0.163 51.47 ;
      END
   END n_4730

   PIN n_8503
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.378 0.163 51.406 ;
      END
   END n_8503

   PIN n_9692
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.978 81.117 13.006 81.28 ;
      END
   END n_9692

   PIN x_out_43_6
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.906 81.117 25.934 81.28 ;
      END
   END x_out_43_6

   PIN FE_OFN130_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.65 81.198 25.678 81.28 ;
      END
   END FE_OFN130_n_27449

   PIN FE_OFN259_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 20.018 81.198 20.046 81.28 ;
      END
   END FE_OFN259_n_4280

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.97 81.198 25.998 81.28 ;
      END
   END ispd_clk

   PIN n_10045
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 28.274 0.163 28.302 ;
      END
   END n_10045

   PIN n_10212
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.186 0.163 51.214 ;
      END
   END n_10212

   PIN n_10216
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.306 0.163 40.334 ;
      END
   END n_10216

   PIN n_10754
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 13.874 0.163 13.902 ;
      END
   END n_10754

   PIN n_11148
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 58.162 0.163 58.19 ;
      END
   END n_11148

   PIN n_12194
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 19.634 0.163 19.662 ;
      END
   END n_12194

   PIN n_12199
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.738 0.163 10.766 ;
      END
   END n_12199

   PIN n_12200
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 62.834 0.163 62.862 ;
      END
   END n_12200

   PIN n_12214
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 40.242 0.163 40.27 ;
      END
   END n_12214

   PIN n_13421
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 45.49 0.163 45.518 ;
      END
   END n_13421

   PIN n_19060
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 54.194 0.163 54.222 ;
      END
   END n_19060

   PIN n_20037
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 23.026 81.117 23.054 81.28 ;
      END
   END n_20037

   PIN n_22693
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.842 81.117 25.87 81.28 ;
      END
   END n_22693

   PIN n_23388
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.898 81.117 22.926 81.28 ;
      END
   END n_23388

   PIN n_24201
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 71.602 0.163 71.63 ;
      END
   END n_24201

   PIN n_24202
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.658 0.163 68.686 ;
      END
   END n_24202

   PIN n_24640
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 68.594 0.163 68.622 ;
      END
   END n_24640

   PIN n_25569
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.906 81.117 25.934 81.28 ;
      END
   END n_25569

   PIN n_26279
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 33.714 81.117 33.742 81.28 ;
      END
   END n_26279

   PIN n_27379
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.482 81.117 34.51 81.28 ;
      END
   END n_27379

   PIN n_27380
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.754 81.117 32.782 81.28 ;
      END
   END n_27380

   PIN n_28713
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.562 81.117 32.59 81.28 ;
      END
   END n_28713

   PIN n_28714
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 32.69 81.117 32.718 81.28 ;
      END
   END n_28714

   PIN n_4859
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.674 0.163 10.702 ;
      END
   END n_4859

   PIN n_6377
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.61 0.163 10.638 ;
      END
   END n_6377

   PIN n_6378
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.546 0.163 10.574 ;
      END
   END n_6378

   PIN n_8054
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.314 0.163 51.342 ;
      END
   END n_8054

   PIN n_8528
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 51.25 0.163 51.278 ;
      END
   END n_8528

   PIN n_8602
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 10.482 0.163 10.51 ;
      END
   END n_8602

   PIN x_in_52_13
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 34.546 81.117 34.574 81.28 ;
      END
   END x_in_52_13

   PIN x_in_52_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 23.026 81.117 23.054 81.28 ;
      END
   END x_in_52_6

   PIN x_out_43_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.594 81.117 28.622 81.28 ;
      END
   END x_out_43_7

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 106.432 81.28 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 106.432 81.28 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 106.432 81.28 ;
      LAYER V1 ;
         RECT 0.0 0.0 106.432 81.28 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 106.432 81.28 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 106.432 81.28 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 106.432 81.28 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 106.432 81.28 ;
      LAYER M1 ;
         RECT 0.0 0.0 106.432 81.28 ;
   END
END h2_mgc_fft_a

MACRO h1_mgc_fft_a
   CLASS BLOCK ;
   FOREIGN h1 ;
   ORIGIN 0 0 ;
   SIZE 97.152 BY 55.04 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1036_n_26168
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 5.362 0.163 5.39 ;
      END
   END FE_OFN1036_n_26168

   PIN n_10017
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 54.642 0.0 54.67 0.163 ;
      END
   END n_10017

   PIN n_11653
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 12.466 54.877 12.494 55.04 ;
      END
   END n_11653

   PIN n_12968
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 37.362 0.0 37.39 0.163 ;
      END
   END n_12968

   PIN n_12983
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.722 0.0 4.75 0.163 ;
      END
   END n_12983

   PIN n_13860
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.706 0.0 54.734 0.163 ;
      END
   END n_13860

   PIN n_14132
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.394 0.0 57.422 0.163 ;
      END
   END n_14132

   PIN n_14219
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 35.058 0.0 35.086 0.163 ;
      END
   END n_14219

   PIN n_14273
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.53 0.0 36.558 0.163 ;
      END
   END n_14273

   PIN n_1985
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.282 0.0 63.31 0.163 ;
      END
   END n_1985

   PIN n_21165
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 89.202 0.0 89.23 0.163 ;
      END
   END n_21165

   PIN n_23487
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.989 30.834 97.152 30.862 ;
      END
   END n_23487

   PIN n_24189
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.802 0.0 74.83 0.163 ;
      END
   END n_24189

   PIN n_24437
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.989 38.962 97.152 38.99 ;
      END
   END n_24437

   PIN n_2458
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.842 0.0 57.87 0.163 ;
      END
   END n_2458

   PIN n_3332
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.522 0.0 57.55 0.163 ;
      END
   END n_3332

   PIN n_4937
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.346 0.0 63.374 0.163 ;
      END
   END n_4937

   PIN n_5596
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 49.586 0.0 49.614 0.163 ;
      END
   END n_5596

   PIN n_5761
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.562 0.0 80.59 0.163 ;
      END
   END n_5761

   PIN n_5771
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.682 0.0 77.71 0.163 ;
      END
   END n_5771

   PIN n_5839
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 57.458 0.0 57.486 0.163 ;
      END
   END n_5839

   PIN n_6223
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 50.546 0.0 50.574 0.163 ;
      END
   END n_6223

   PIN n_6579
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.986 0.0 40.014 0.163 ;
      END
   END n_6579

   PIN n_6722
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 69.042 0.0 69.07 0.163 ;
      END
   END n_6722

   PIN n_7868
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.674 0.0 74.702 0.163 ;
      END
   END n_7868

   PIN n_7889
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 48.882 0.0 48.91 0.163 ;
      END
   END n_7889

   PIN n_8086
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 17.266 0.0 17.294 0.163 ;
      END
   END n_8086

   PIN n_8089
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.706 0.0 62.734 0.163 ;
      END
   END n_8089

   PIN n_8142
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 46.002 0.0 46.03 0.163 ;
      END
   END n_8142

   PIN n_8523
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 71.922 0.0 71.95 0.163 ;
      END
   END n_8523

   PIN n_8596
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.186 0.0 43.214 0.163 ;
      END
   END n_8596

   PIN n_8597
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 43.122 0.0 43.15 0.163 ;
      END
   END n_8597

   PIN n_8601
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.762 0.0 51.79 0.163 ;
      END
   END n_8601

   PIN n_8972
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.602 0.0 31.63 0.163 ;
      END
   END n_8972

   PIN x_out_29_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.989 22.322 97.152 22.35 ;
      END
   END x_out_29_0

   PIN x_out_29_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.882 0.163 16.91 ;
      END
   END x_out_29_1

   PIN x_out_37_21
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.989 28.018 97.152 28.046 ;
      END
   END x_out_37_21

   PIN x_out_38_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.989 30.834 97.152 30.862 ;
      END
   END x_out_38_12

   PIN x_out_6_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.989 36.594 97.152 36.622 ;
      END
   END x_out_6_10

   PIN x_out_6_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.989 19.314 97.152 19.342 ;
      END
   END x_out_6_11

   PIN FE_OFN251_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 22.002 54.958 22.03 55.04 ;
      END
   END FE_OFN251_n_4162

   PIN FE_OFN306_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.282 0.082 39.31 ;
      END
   END FE_OFN306_n_3069

   PIN FE_OFN324_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 97.07 39.282 97.152 39.31 ;
      END
   END FE_OFN324_n_4860

   PIN FE_OFN330_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 74.802 54.958 74.83 55.04 ;
      END
   END FE_OFN330_n_4860

   PIN FE_OFN393_n_14663
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 16.946 54.877 16.974 55.04 ;
      END
   END FE_OFN393_n_14663

   PIN FE_OFN662_n_27899
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.65 0.163 49.678 ;
      END
   END FE_OFN662_n_27899

   PIN FE_OFN810_n_12878
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.989 16.562 97.152 16.59 ;
      END
   END FE_OFN810_n_12878

   PIN FE_OFN93_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 16.626 0.082 16.654 ;
      END
   END FE_OFN93_n_27449

   PIN FE_OFN96_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.33 0.082 49.358 ;
      END
   END FE_OFN96_n_27449

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.25 0.082 27.278 ;
      END
   END ispd_clk

   PIN n_10004
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 72.498 0.0 72.526 0.163 ;
      END
   END n_10004

   PIN n_12575
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 59.762 0.0 59.79 0.163 ;
      END
   END n_12575

   PIN n_13218
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.802 0.0 74.83 0.163 ;
      END
   END n_13218

   PIN n_13671
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.034 0.0 74.062 0.163 ;
      END
   END n_13671

   PIN n_13859
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.642 0.0 54.67 0.163 ;
      END
   END n_13859

   PIN n_14448
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.738 0.0 74.766 0.163 ;
      END
   END n_14448

   PIN n_14791
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.642 0.0 70.67 0.163 ;
      END
   END n_14791

   PIN n_17925
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 4.658 54.877 4.686 55.04 ;
      END
   END n_17925

   PIN n_21076
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 97.07 13.554 97.152 13.582 ;
      END
   END n_21076

   PIN n_21393
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.09 0.163 39.118 ;
      END
   END n_21393

   PIN n_21394
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 39.026 0.163 39.054 ;
      END
   END n_21394

   PIN n_21551
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 84.466 0.0 84.494 0.163 ;
      END
   END n_21551

   PIN n_23020
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 9.842 54.877 9.87 55.04 ;
      END
   END n_23020

   PIN n_2355
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 60.402 0.0 60.43 0.163 ;
      END
   END n_2355

   PIN n_24577
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 38.962 0.163 38.99 ;
      END
   END n_24577

   PIN n_25555
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 36.594 0.163 36.622 ;
      END
   END n_25555

   PIN n_25843
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 27.122 0.163 27.15 ;
      END
   END n_25843

   PIN n_26168
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 96.989 3.122 97.152 3.15 ;
      END
   END n_26168

   PIN n_26689
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 34.482 0.163 34.51 ;
      END
   END n_26689

   PIN n_28608
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 49.458 0.082 49.486 ;
      END
   END n_28608

   PIN n_2901
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 66.418 0.0 66.446 0.163 ;
      END
   END n_2901

   PIN n_4914
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.578 0.0 54.606 0.163 ;
      END
   END n_4914

   PIN n_5242
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 72.882 0.0 72.91 0.163 ;
      END
   END n_5242

   PIN n_5597
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 80.626 0.0 80.654 0.163 ;
      END
   END n_5597

   PIN n_5828
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 56.242 0.0 56.27 0.163 ;
      END
   END n_5828

   PIN n_7867
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.682 0.0 77.71 0.163 ;
      END
   END n_7867

   PIN n_8074
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 70.322 0.0 70.35 0.163 ;
      END
   END n_8074

   PIN n_8076
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.858 0.0 71.886 0.163 ;
      END
   END n_8076

   PIN n_8650
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 63.218 0.0 63.246 0.163 ;
      END
   END n_8650

   PIN n_8971
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 31.346 0.0 31.374 0.163 ;
      END
   END n_8971

   PIN n_9998
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 74.866 0.0 74.894 0.163 ;
      END
   END n_9998

   PIN n_9999
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.746 0.0 77.774 0.163 ;
      END
   END n_9999

   PIN x_in_46_0
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 96.989 22.258 97.152 22.286 ;
      END
   END x_in_46_0

   PIN x_in_61_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 48.882 0.0 48.91 0.082 ;
      END
   END x_in_61_5

   PIN x_in_61_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 43.314 0.0 43.342 0.082 ;
      END
   END x_in_61_6

   PIN x_in_61_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 59.698 0.0 59.726 0.082 ;
      END
   END x_in_61_7

   PIN x_in_61_8
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 66.61 0.0 66.638 0.082 ;
      END
   END x_in_61_8

   PIN x_in_61_9
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 69.042 0.0 69.07 0.082 ;
      END
   END x_in_61_9

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 97.152 55.04 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 97.152 55.04 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 97.152 55.04 ;
      LAYER V1 ;
         RECT 0.0 0.0 97.152 55.04 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 97.152 55.04 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 97.152 55.04 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 97.152 55.04 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 97.152 55.04 ;
      LAYER M1 ;
         RECT 0.0 0.0 97.152 55.04 ;
   END
END h1_mgc_fft_a

MACRO h0_mgc_fft_a
   CLASS BLOCK ;
   FOREIGN h0 ;
   ORIGIN 0 0 ;
   SIZE 105.472 BY 50.56 ;
   SYMMETRY X Y R90 ;
   PIN n_13301
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 54.962 0.0 54.99 0.163 ;
      END
   END n_13301

   PIN n_13302
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.122 0.0 51.15 0.163 ;
      END
   END n_13302

   PIN n_13303
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 51.186 0.0 51.214 0.163 ;
      END
   END n_13303

   PIN n_13488
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 71.346 0.0 71.374 0.163 ;
      END
   END n_13488

   PIN n_14077
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 79.282 0.0 79.31 0.163 ;
      END
   END n_14077

   PIN n_14078
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.106 0.0 77.134 0.163 ;
      END
   END n_14078

   PIN n_14581
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 77.106 0.0 77.134 0.163 ;
      END
   END n_14581

   PIN n_15640
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 39.666 0.0 39.694 0.163 ;
      END
   END n_15640

   PIN n_15661
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 68.466 0.0 68.494 0.163 ;
      END
   END n_15661

   PIN n_16544
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.618 0.0 77.646 0.163 ;
      END
   END n_16544

   PIN n_19438
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 105.309 7.218 105.472 7.246 ;
      END
   END n_19438

   PIN n_20533
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 105.309 25.586 105.472 25.614 ;
      END
   END n_20533

   PIN n_3465
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.97 0.0 17.998 0.163 ;
      END
   END n_3465

   PIN n_6033
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.386 0.0 30.414 0.163 ;
      END
   END n_6033

   PIN n_7083
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.266 0.0 25.294 0.163 ;
      END
   END n_7083

   PIN n_7084
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.33 0.0 25.358 0.163 ;
      END
   END n_7084

   PIN x_out_15_20
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 61.234 50.397 61.262 50.56 ;
      END
   END x_out_15_20

   PIN x_out_15_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 105.309 41.01 105.472 41.038 ;
      END
   END x_out_15_24

   PIN FE_OFN1111_rst
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 105.39 8.946 105.472 8.974 ;
      END
   END FE_OFN1111_rst

   PIN FE_OFN17_n_29617
      DIRECTION INPUT ;
      PORT 
         LAYER MINT3 ;
             RECT 0.0 8.818 0.163 8.846 ;
      END
   END FE_OFN17_n_29617

   PIN FE_OFN251_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.21 0.0 100.238 0.082 ;
      END
   END FE_OFN251_n_4162

   PIN FE_OFN288_n_29266
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 86.578 0.0 86.606 0.163 ;
      END
   END FE_OFN288_n_29266

   PIN FE_OFN314_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 76.978 0.0 77.006 0.082 ;
      END
   END FE_OFN314_n_3069

   PIN FE_OFN409_n_28303
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 0.0 43.89 0.082 43.918 ;
      END
   END FE_OFN409_n_28303

   PIN FE_OFN660_n_19445
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 88.626 0.0 88.654 0.163 ;
      END
   END FE_OFN660_n_19445

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 42.866 0.0 42.894 0.082 ;
      END
   END ispd_clk

   PIN n_10314
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 30.962 0.0 30.99 0.163 ;
      END
   END n_10314

   PIN n_10315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 36.786 0.0 36.814 0.163 ;
      END
   END n_10315

   PIN n_11856
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 85.362 0.0 85.39 0.163 ;
      END
   END n_11856

   PIN n_15273
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 62.706 0.0 62.734 0.163 ;
      END
   END n_15273

   PIN n_17533
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 100.082 0.0 100.11 0.163 ;
      END
   END n_17533

   PIN n_18413
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 77.042 0.0 77.07 0.163 ;
      END
   END n_18413

   PIN n_20363
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 100.082 0.0 100.11 0.163 ;
      END
   END n_20363

   PIN n_21988
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 103.73 0.0 103.758 0.082 ;
      END
   END n_21988

   PIN n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 105.39 25.458 105.472 25.486 ;
      END
   END n_27449

   PIN n_3028
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 17.906 0.0 17.934 0.163 ;
      END
   END n_3028

   PIN n_3132
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.29 0.0 18.318 0.163 ;
      END
   END n_3132

   PIN n_3771
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 28.082 0.0 28.11 0.163 ;
      END
   END n_3771

   PIN n_4593
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.194 0.0 22.222 0.163 ;
      END
   END n_4593

   PIN n_4594
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.002 0.0 22.03 0.163 ;
      END
   END n_4594

   PIN n_4873
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 19.442 0.0 19.47 0.163 ;
      END
   END n_4873

   PIN n_5057
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 22.258 0.0 22.286 0.163 ;
      END
   END n_5057

   PIN n_5315
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 18.162 0.0 18.19 0.163 ;
      END
   END n_5315

   PIN n_6966
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 25.202 0.0 25.23 0.163 ;
      END
   END n_6966

   PIN n_7082
      DIRECTION INPUT ;
      PORT 
         LAYER MINT2 ;
             RECT 27.378 0.0 27.406 0.163 ;
      END
   END n_7082

   PIN n_871
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 105.309 8.818 105.472 8.846 ;
      END
   END n_871

   PIN x_in_25_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 25.202 0.0 25.23 0.082 ;
      END
   END x_in_25_4

   PIN x_in_25_5
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 18.098 0.0 18.126 0.082 ;
      END
   END x_in_25_5

   PIN x_in_25_6
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 30.77 0.0 30.798 0.082 ;
      END
   END x_in_25_6

   PIN x_in_25_7
      DIRECTION INPUT ;
      PORT 
         LAYER MINT4 ;
             RECT 3.058 0.0 3.086 0.082 ;
      END
   END x_in_25_7

   PIN x_out_38_4
      DIRECTION INPUT ;
      PORT 
         LAYER MINT1 ;
             RECT 105.309 20.85 105.472 20.878 ;
      END
   END x_out_38_4

   OBS
      LAYER VINT3 ;
         RECT 0.0 0.0 105.472 50.56 ;
      LAYER VINT2 ;
         RECT 0.0 0.0 105.472 50.56 ;
      LAYER VINT1 ;
         RECT 0.0 0.0 105.472 50.56 ;
      LAYER V1 ;
         RECT 0.0 0.0 105.472 50.56 ;
      LAYER MINT4 ;
         RECT 0.0 0.0 105.472 50.56 ;
      LAYER MINT3 ;
         RECT 0.0 0.0 105.472 50.56 ;
      LAYER MINT2 ;
         RECT 0.0 0.0 105.472 50.56 ;
      LAYER MINT1 ;
         RECT 0.0 0.0 105.472 50.56 ;
      LAYER M1 ;
         RECT 0.0 0.0 105.472 50.56 ;
   END
END h0_mgc_fft_a

END LIBRARY 
